`timescale 1ns / 1ps

module tb;

    parameter SYS_PERIOD = 10;    //clk 100M, 10ns (fixed)
    
    reg clk, rst;
    reg [127:0] state, key;
    wire [127:0] out;
    
    //clock generation (fixed)
    initial begin
        forever
        #(SYS_PERIOD/2) clk = ~clk;
    end
    
    aes_top DUT (.clk(clk), .state(state), .key(key), .out(out), .rst(rst));
    
    initial begin
        clk = 0;
        rst = 0;
        #10
        rst = 1;
        #10
        rst = 0;
        key = 128'hcd32_fe58_4188_9413_8499_ef35_6910_c98d;
        state = 128'h296d_e070_6aa6_af23_1ecb_3dbe_f494_bc16;

        #200;
        key = 128'h2111_382d_46a7_f295_747d_6616_ea48_02f1;
        state = 128'hd8ed_651c_91b1_649a_5533_c9eb_7ae9_6a15;

        #200;
        key = 128'h1544_526b_e7fb_6717_448f_09c2_483f_26eb;
        state = 128'h7682_334c_d4ac_62e5_33e5_2569_cb5a_e4d7;

        #200;
        key = 128'h0f1c_0d59_d70c_ec84_75aa_e83f_f57f_650f;
        state = 128'h6e84_22ff_417b_8bd5_3f94_e79d_bfe2_3b10;

        #200;
        key = 128'hf03a_340d_890a_dc71_b47a_eebd_5606_bf88;
        state = 128'h4975_97d1_0afd_95cf_c4f1_620e_e75d_5b87;

        #200;
        key = 128'hc222_c62f_915d_3b21_dbbc_75ff_e117_2b5b;
        state = 128'h8515_fdab_31fd_b21e_666a_799b_8b1e_eca6;

        #200;
        key = 128'h8d49_9f8b_f9f9_9f27_c8d7_7d59_d014_8c06;
        state = 128'h973c_dfa6_f46b_36af_12d4_bebe_9343_16b1;

        #200;
        key = 128'h7d28_eba7_a699_aa23_6db6_b18b_cafe_f82f;
        state = 128'h7f02_82e1_9ebb_3551_dc65_5b96_e2ff_df98;

        #200;
        key = 128'he3b4_d673_4d29_bf1c_dc9f_1d8b_44d9_59b6;
        state = 128'h6987_0951_ad5d_2de0_2b96_3255_6118_0f6f;

        #200;
        key = 128'h6edf_bc2f_c3de_bc8e_4941_c649_793a_9c0f;
        state = 128'h3962_04d6_f4db_4d17_5382_6e5c_78e7_d198;

        #200;
        key = 128'h2681_1316_9f45_a87b_f347_f1dc_aebb_8263;
        state = 128'h492d_6e64_8cbd_e23e_e49b_e20d_e077_361d;

        #200;
        key = 128'hb7dc_c22e_8336_24d7_a22f_f906_c309_db44;
        state = 128'h522c_41b0_f441_75c0_c554_8754_9fc7_4238;

        #200;
        key = 128'hf4b9_c291_74b0_0a10_8b4b_42ff_a45b_61e1;
        state = 128'h23c2_c757_2765_7835_3593_241f_c655_a050;

        #200;
        key = 128'hd541_11b4_45d2_9785_bd9a_40ba_629e_7b88;
        state = 128'h1ba9_c87b_912a_fbaa_c96b_08fc_2da5_471f;

        #200;
        key = 128'h5783_143a_2478_dde6_1396_c578_3daa_679c;
        state = 128'hd08d_eb74_9bca_86a6_57e5_ee0f_189f_7543;

        #200;
        key = 128'h1dc2_9ffd_a463_e5e0_ed20_8443_0421_283d;
        state = 128'h4fa2_68d5_96ab_fb21_55d1_eac7_464e_5094;

        #200;
        key = 128'h5c11_711d_f9e5_efcc_8b40_c9d1_b5a2_0848;
        state = 128'h0a20_3b1a_cb31_8c3d_b3ea_dc07_2c51_a832;

        #200;
        key = 128'h0e3a_52f6_66fc_b412_5a26_2c2d_8e6c_a00e;
        state = 128'h311c_7d2e_a59b_c53c_65c1_462f_dff4_c65c;

        #200;
        key = 128'h5923_e82f_e9cc_aaf5_1611_5482_57a8_5a06;
        state = 128'h24d6_1007_1c6d_3e5e_2e4e_27d6_26d2_256c;

        #200;
        key = 128'h4b67_2c98_b1a7_a15d_3ba7_6af2_90a4_f342;
        state = 128'h5ade_6db3_da19_d752_11ad_0fa2_c563_ffd2;

        #200;
        key = 128'h4cf7_1904_84ae_fbcd_cf08_bb3a_6fd5_a152;
        state = 128'hdee5_e9bc_cad3_7763_4ee6_8491_40d9_c129;

        #200;
        key = 128'h1024_0051_ea88_9297_8cf3_b77e_df63_3d70;
        state = 128'h2eec_86d9_61b2_c285_f260_9110_ae2b_3d86;

        #200;
        key = 128'h0578_99b9_261e_0010_f345_8f72_04d6_a508;
        state = 128'ha4c1_e91f_190b_fc9e_6190_80d8_a166_7289;

        #200;
        key = 128'he0f7_cef0_25f3_81d2_b7d1_f4e4_d617_8472;
        state = 128'h502a_ca6b_4bfd_a62b_0365_631c_04fc_eaa1;

        #200;
        key = 128'h5b27_027b_0b3e_9f41_2bc6_a2c2_cbab_e816;
        state = 128'h5573_fe81_9d08_7d50_6fc7_6ade_ec44_799e;

        #200;
        key = 128'he37c_a8e1_0e7f_51a9_8b48_88d2_6ce4_0418;
        state = 128'h8710_a1fe_54d5_6688_308d_b31b_25f6_10e4;

        #200;
        key = 128'h3db3_8693_1ae6_c36b_596f_6383_e6d0_e3c0;
        state = 128'h8661_8b12_cbb3_6dc0_bca5_9320_9edb_181e;

        #200;
        key = 128'hf611_415e_3257_ce98_baa8_73e1_4fd4_bf39;
        state = 128'h905b_726c_e830_a8aa_8429_493c_5cd6_ec8c;

        #200;
        key = 128'h4420_cf7f_fe88_77fe_8726_ac55_8d10_bf3a;
        state = 128'hd2be_f96c_5f68_a420_4320_2de8_f7e9_1b2b;

        #200;
        key = 128'hbf79_a718_1e81_f1de_ea1d_4681_232d_9e07;
        state = 128'hf392_7605_a262_b981_4fc1_a927_bea8_f840;

        #200;
        key = 128'hfcd4_d409_965c_6068_5eae_2edc_0933_3e72;
        state = 128'h9576_e1a2_ef6a_dae6_21db_cd80_a000_b8b6;

        #200;
        key = 128'h9411_d9b9_65cd_273a_e2ee_f4f8_c531_046a;
        state = 128'hc597_5274_a3bd_adfc_00d5_8404_4294_ea28;

        #200;
        key = 128'hc2b0_ed12_130c_0a14_2433_ef16_c737_f5d0;
        state = 128'ha499_a121_81e6_25a8_2b2b_e086_ec24_d473;

        #200;
        key = 128'h423c_05b1_2ba8_fd3b_d9ad_d358_821b_c532;
        state = 128'h7e68_09c3_bfb0_ebec_4da5_b15a_1ece_12d3;

        #200;
        key = 128'h3e68_57bd_582e_8a1f_89c6_6622_b645_5876;
        state = 128'hf89e_98f1_7302_6be2_690f_c692_3947_03b6;

        #200;
        key = 128'h5a57_5d94_a1a5_d314_c5f9_ffbb_35af_ab3e;
        state = 128'h42ea_9873_d3c5_4055_0878_f6c8_289c_aac4;

        #200;
        key = 128'h7a2b_8355_af56_ff26_4964_e2ac_05b9_1167;
        state = 128'h824d_59e7_8db9_96e9_051d_c64e_cfbb_dac7;

        #200;
        key = 128'h62bb_5cae_8d54_2bd6_8e9b_6cc5_9e2a_a83c;
        state = 128'hc1a4_44fb_fa55_ef2f_7a21_1a6d_8f6e_35d6;

        #200;
        key = 128'h5796_c4b3_d22d_d766_ee4c_798d_3667_5abb;
        state = 128'h6b31_2635_08e0_4636_3798_9a55_ea5e_109a;

        #200;
        key = 128'h58f7_eb9d_2d74_80d8_1fc8_22d6_64c6_c719;
        state = 128'hbd49_af52_8245_bfed_cb1b_9ee6_5f3c_28a8;

        #200;
        key = 128'h7e2b_9bd5_2227_7ec0_024e_820f_8be1_82ab;
        state = 128'hf9ba_6b82_09d1_b84d_f111_ed51_1dd3_c0ef;

        #200;
        key = 128'h976e_1782_f7ab_55b5_fd23_e7a3_8db5_c6c0;
        state = 128'h39c2_f92a_daef_81f4_58c4_7ff4_190e_baaf;

        #200;
        key = 128'h8758_1a3a_ed10_4ff4_8f3b_1419_9748_9edb;
        state = 128'hd983_d0ce_ddf0_b160_cfb6_3890_e2b3_046c;

        #200;
        key = 128'h1a0d_4603_7554_f5f6_556a_cdac_ec12_997a;
        state = 128'h030f_d648_4337_046e_8e53_e0ea_df32_8711;

        #200;
        key = 128'h5cd5_a02f_14c4_e3e4_d4cb_45c6_e690_da9b;
        state = 128'h9fbe_9a4d_9d63_573e_cf1f_8998_3232_7c95;

        #200;
        key = 128'h2a6c_2d36_b8f9_d065_445f_92ed_5503_497e;
        state = 128'hef36_a61a_fc57_8b91_98c7_b971_a326_b2ce;

        #200;
        key = 128'h7b39_3edd_e46e_3987_dede_0351_796f_f6f8;
        state = 128'h9378_6122_b5ae_e2df_2b20_30e5_3ebd_2c6e;

        #200;
        key = 128'heb97_190b_261c_bb50_ffea_61a0_4d22_da9a;
        state = 128'h2b0b_0891_639e_f0ff_2b54_e08e_4cae_7fc8;

        #200;
        key = 128'h85d9_3c04_e34f_c585_2248_4e27_e8bc_275b;
        state = 128'h43b9_9bd7_263a_9da1_e07f_b5af_0f37_d122;

        #200;
        key = 128'h0dd2_6cfe_3f8a_84d1_d572_1f17_8b3c_890f;
        state = 128'hb452_02a5_1088_b3fe_6118_c16d_1799_87db;

        #200;
        key = 128'h81ee_7a72_7614_da91_7636_da76_61c6_5da0;
        state = 128'h8171_4a78_638e_86d9_900c_c882_d6d5_01eb;

        #200;
        key = 128'hdfb8_74c7_c393_fa53_4954_2344_9256_14c9;
        state = 128'h8f3d_be49_2400_1695_ad7f_3f17_874e_9497;

        #200;
        key = 128'ha485_8222_b416_f4ab_d46e_0944_db1d_e154;
        state = 128'heb30_4610_e5ac_617d_8494_c03b_119a_8131;

        #200;
        key = 128'h2eb7_080c_66b3_a467_5c53_298f_e13a_7a5b;
        state = 128'haf7d_b321_3363_6bc0_f58a_ff4a_f4a2_1e23;

        #200;
        key = 128'h8b62_ed4d_deb6_04ee_a918_9221_942f_fbdf;
        state = 128'h64e0_80d5_3981_5456_1677_fc81_1e4d_f526;

        #200;
        key = 128'hc5dc_71de_b794_2990_6933_55df_312f_145d;
        state = 128'h4062_8548_28d5_8b6a_461c_38fb_1c50_4e8d;

        #200;
        key = 128'h5fb4_1d12_9226_30e1_2456_9487_f787_68a8;
        state = 128'h1c1a_404d_7355_0f9f_90fe_9c37_cfef_2b91;

        #200;
        key = 128'h6585_da70_7d3f_6c8a_8ea6_0d50_5834_519d;
        state = 128'hbdb5_10ae_f9b7_19d9_c77f_0fb1_d491_6c85;

        #200;
        key = 128'h9223_342d_eed5_9e41_2de1_f5c6_7c5a_7508;
        state = 128'h3696_31f0_3123_9d80_e605_12c1_3e06_60c1;

        #200;
        key = 128'he3bd_cbb6_7f2b_cf90_907b_8d9f_ff70_98a8;
        state = 128'h770b_a291_ec0b_1b5c_ca0b_2313_88ca_e9ed;

        #200;
        key = 128'ha1e3_5d8c_c6a8_9565_e55b_6c87_d26a_42ca;
        state = 128'h6e3f_e701_4f0e_8414_8e3e_6844_eef1_26ad;

        #200;
        key = 128'h866f_9bbc_422a_7913_7a90_3c10_1fcc_6ac6;
        state = 128'h45d3_8073_736c_1d1a_e265_3051_fa01_afd7;

        #200;
        key = 128'h9d8f_7128_c01c_e972_5cfc_2629_bc31_e0df;
        state = 128'h9862_dddf_6f10_0f39_b737_3722_fa3e_34da;

        #200;
        key = 128'ha330_a08f_9d7e_37ad_e147_9d6b_be9e_c784;
        state = 128'haeff_2ff2_dbbf_84e3_f882_7acc_f0df_9fbe;

        #200;
        key = 128'h8053_a220_1d99_a5c8_4e1a_ee01_b2e6_ee61;
        state = 128'hbcbd_3bdd_da98_d0d4_c92e_a555_f61e_3c13;

        #200;
        key = 128'h7211_89c4_5e33_966e_507e_b0ec_d35c_2b94;
        state = 128'ha90a_0156_8efe_5c8b_da33_3408_02e3_4ead;

        #200;
        key = 128'hf96b_7476_6250_32c1_a1c1_3eda_3730_7858;
        state = 128'hd857_35c6_e949_7868_a9fb_5831_b5dd_c891;

        #200;
        key = 128'hd20f_63e1_5609_5fa3_c2ca_a6ba_f6ac_9ea1;
        state = 128'h659e_0a58_a94a_1db9_7157_385b_3f20_d2af;

        #200;
        key = 128'h6747_b263_a031_d4e8_54c0_4aa1_1c73_9994;
        state = 128'h06a7_6a67_2055_00c4_6bca_f81b_9544_37e9;

        #200;
        key = 128'h1c0b_c53b_1788_d7dd_f2f8_17b8_cf8a_4cbf;
        state = 128'h6e38_62c2_642f_49a7_a0d1_11d3_d5eb_8bd3;

        #200;
        key = 128'hcccf_25c2_df0d_a18c_34c3_3a36_1390_0195;
        state = 128'h7599_5bad_5c10_e8c6_1e5a_2a59_d37d_7a4f;

        #200;
        key = 128'h410b_4d41_78a2_47fc_d38f_d2ce_f295_57f9;
        state = 128'he21c_1001_ebe1_0d37_fd0b_b429_6b98_518a;

        #200;
        key = 128'ha91d_6d5d_7da8_0bb6_4f09_ab5b_2b20_55dd;
        state = 128'h3711_3923_2c56_0726_3efa_a52f_b137_b18f;

        #200;
        key = 128'he471_07ed_1a7a_4e6b_39dc_b597_15c7_4e18;
        state = 128'h9b61_9f69_fd83_8dbc_d5e1_8e81_c893_282a;

        #200;
        key = 128'h04f5_2567_6401_ea74_fc6b_860a_93c5_4395;
        state = 128'h989d_147f_56ee_6640_c8d4_a3de_dede_4786;

        #200;
        key = 128'h7ec0_d627_e085_cb19_0efb_47dc_765d_29d1;
        state = 128'h4a54_0021_53b0_24cf_1a69_f0cc_ed14_03b7;

        #200;
        key = 128'h122f_b7ec_c1c0_34c8_a197_a50d_d24a_4350;
        state = 128'h4a2e_0cf0_3c50_3bbc_e1f7_a25b_f1ce_87f3;

        #200;
        key = 128'h6c5c_0b39_4205_9434_fc40_72f3_6da6_6018;
        state = 128'h9d3c_8d00_bdcf_2cf9_c8c7_7673_d550_7be2;

        #200;
        key = 128'h3946_ed19_782c_8b41_f7e8_d2e7_37ed_276a;
        state = 128'hd7c0_e7b0_54fc_725e_8496_2369_5568_c453;

        #200;
        key = 128'hfdfd_b372_c326_7974_9e92_d154_032d_aeae;
        state = 128'ha437_97f6_c330_60d8_ba3f_13ba_ad65_e9bd;

        #200;
        key = 128'h9fd7_f6bf_093c_5d56_03bd_b448_3b7c_8087;
        state = 128'h584e_b253_abbe_378e_dc84_aa56_a66b_a36f;

        #200;
        key = 128'h55b5_33df_187e_99b0_8c26_91f4_6825_ac44;
        state = 128'hba2a_5c4d_6181_d918_7aa6_8824_64af_2f19;

        #200;
        key = 128'h3e79_d18c_d8cd_32cf_eb14_5d5a_5484_155c;
        state = 128'hf94b_eb86_64ad_5b64_723f_539e_2382_4520;

        #200;
        key = 128'h5955_ca90_993d_33b4_df3d_25aa_b3f0_9a70;
        state = 128'h941c_49ce_da3b_df45_b80d_2445_7b25_f53a;

        #200;
        key = 128'hdcb5_99c3_95f7_d383_649e_d27a_7a0d_973d;
        state = 128'h4c82_213b_2d55_7713_8c8a_4d35_733d_679d;

        #200;
        key = 128'h5eb1_ca93_a38d_fdfa_70a5_437b_be9f_b783;
        state = 128'h4921_b66d_b0c4_9aa9_6f28_2a80_a9e8_7752;

        #200;
        key = 128'h1f95_aa3c_926b_a4f0_6a08_b37d_0b57_93d3;
        state = 128'h45cf_b2de_6064_78fa_2a27_1627_b98f_9afb;

        #200;
        key = 128'h666c_2b5a_47dc_5a38_9d71_0d42_0a1d_9bcb;
        state = 128'h40f1_ec64_b3e1_c06c_b20c_19b6_753a_4ac6;

        #200;
        key = 128'hdf9c_a843_8201_2848_c832_9da0_4433_1b3b;
        state = 128'hcfad_db13_31b7_8216_9331_12cf_52f6_19a8;

        #200;
        key = 128'h9417_b9fb_8e9d_5251_0280_a1e4_3a77_6212;
        state = 128'hc4e4_7c9f_0ad9_d4af_9fdd_b775_65ef_3632;

        #200;
        key = 128'hf1b1_f468_c5c7_b319_2baf_be53_a25a_fbf4;
        state = 128'hec11_35a1_295a_a91b_36da_5bda_10e6_ecbc;

        #200;
        key = 128'he63c_1ddf_cc21_8bac_e56f_852b_4bb9_07d9;
        state = 128'h4282_ac43_9fab_5dd8_33a6_1d33_9298_29ae;

        #200;
        key = 128'hb1f9_6c2f_3031_71c6_f1d1_7c2d_b1c0_0ac7;
        state = 128'h5c0b_7332_afaf_7657_8edd_e3f7_ef0e_ce28;

        #200;
        key = 128'h27a2_9f51_7e4d_24b4_47b5_7d22_3a70_e0a0;
        state = 128'h02ac_efd2_dc4f_4d3b_30ed_c767_12ab_b1bd;

        #200;
        key = 128'h7584_690b_6afd_6f7e_55ad_123a_3a61_189d;
        state = 128'h7a01_a646_200f_8ef1_591a_634c_6919_e7b8;

        #200;
        key = 128'h9f7e_12b8_b995_5b2d_be9b_5a03_d69b_580f;
        state = 128'h2d32_fee9_3699_3958_b1eb_14a0_bd23_4c8a;

        #200;
        key = 128'h0181_4818_dce9_06c7_2d19_2ac9_f88f_7261;
        state = 128'hcabf_5144_fd38_2057_4b0f_d2a4_b8f9_0e69;

        #200;
        key = 128'h5e05_f421_4add_079e_71f5_668e_9464_9a8c;
        state = 128'h1e7a_f14b_b2cf_47e4_4b04_1db0_40ca_0ce6;

        #200;
        key = 128'heceb_c1e8_0cb3_a06a_0c7b_8c1a_e4ba_77aa;
        state = 128'h0369_2389_6713_d2c9_a7aa_7782_5aa9_25c4;

        #200;
        key = 128'h09ad_e01a_0a8d_b545_8b00_55c2_acd2_566e;
        state = 128'hf41a_40bc_3f59_83ca_7a13_2e18_6196_bf7b;

        #200;
        key = 128'h4228_ff9a_5e44_8d6f_3299_65f5_3ac1_0124;
        state = 128'hf4ce_1941_5c20_c3dd_6103_8571_53d7_9bc2;

        #200;
        key = 128'hd264_e327_1aa8_c2ef_89d1_9d4e_1fa3_8b68;
        state = 128'h6245_e681_a9fb_a837_7bef_05d4_eb63_ddf2;

        #200;
        key = 128'ha443_ebf6_0fdb_6e2c_5df4_7157_e0e5_4ea4;
        state = 128'h43ad_c402_e29f_9d05_80e3_7378_00ed_d56c;

        #200;
        key = 128'h54f3_c99f_90f3_a563_acd0_06ba_38df_20a9;
        state = 128'h001d_0578_96a8_94eb_ef57_d38c_b189_45dd;

        #200;
        key = 128'h3410_15da_c0c9_c4ae_fcbd_3a52_6c00_5f1f;
        state = 128'ha1bf_5936_eb99_fe83_8f41_bb97_27ad_463f;

        #200;
        key = 128'h9270_e16d_d20e_9b02_cf4c_9d44_1a9d_f7ef;
        state = 128'h5616_f269_219b_8c83_9ea8_fd70_6738_5bd0;

        #200;
        key = 128'he5eb_37ac_8741_0fc9_701b_5570_4a9f_6688;
        state = 128'h7256_8360_c38d_1888_42c9_55ba_1c15_9144;

        #200;
        key = 128'h111b_dd7c_3645_66dc_1dd6_0ad4_7f1d_1e5d;
        state = 128'h57d3_9608_f52c_54f3_7605_7a9b_d409_d5e8;

        #200;
        key = 128'h8e5b_55ff_15bd_7a8c_a544_abcc_7dc0_04ae;
        state = 128'h0cc4_05b5_c2db_5506_6602_df9c_e193_bfc5;

        #200;
        key = 128'h486b_8942_563c_ddb5_b3cd_fb6f_6fa8_be47;
        state = 128'hadbc_0d51_18ef_623f_8f3e_a93c_8403_8862;

        #200;
        key = 128'ha353_339c_c574_16a6_3f16_b129_c684_f4fa;
        state = 128'h1d6c_2ad8_7c98_b519_2c79_2f1f_cc79_c11d;

        #200;
        key = 128'hcb5b_02dd_ee16_7168_0878_e58f_8ffd_f43b;
        state = 128'h59e9_0644_8c08_95ae_c034_f9ad_c891_db49;

        #200;
        key = 128'he02d_208b_4d5c_aef6_b6c0_1f3c_8c6d_bea3;
        state = 128'h601d_1160_f37f_db84_fd0e_3c5b_a61b_e97b;

        #200;
        key = 128'h318b_3323_9c84_66ad_b063_8027_bb5a_ab72;
        state = 128'h36ce_56c7_4361_1c80_651e_bd49_8687_4ba6;

        #200;
        key = 128'hf20c_2c74_1cf4_db55_0e8d_0f2b_a1c9_a3da;
        state = 128'h3f58_ecc6_da22_c3c8_8b70_8131_58d4_7060;

        #200;
        key = 128'he1f8_4591_a622_f5ee_dc7f_a8c7_2cd3_c044;
        state = 128'hab10_b467_e70f_ef0e_a0cf_1937_1473_23cb;

        #200;
        key = 128'hace0_d72f_0aa5_c302_129c_b136_5876_b7e3;
        state = 128'h7da9_af2b_20a1_8e29_dc6c_fc52_d264_7ed5;

        #200;
        key = 128'h007b_7e82_e489_6344_f64b_b188_8a25_034c;
        state = 128'ha45d_1bb4_e806_8801_4656_dc5d_fda8_dc1b;

        #200;
        key = 128'h7b4e_08da_7ef2_e3e5_09cf_2c48_2297_5cad;
        state = 128'h1a45_a8b3_70d4_f45f_2113_af19_b1c1_0490;

        #200;
        key = 128'hd2e6_fa5b_9833_eb5c_41bf_a489_dce5_f413;
        state = 128'hcd51_3f1f_92e1_ee65_2aac_a149_4f52_9ae5;

        #200;
        key = 128'h9c06_07b2_07cc_334d_8515_6c14_394f_a3b2;
        state = 128'hd2ff_f293_e7e3_d6cc_4ae5_d74b_1e40_2920;

        #200;
        key = 128'h4f50_d320_f810_448b_cbac_7b2a_95c1_de0e;
        state = 128'h0140_de40_fc90_663d_719d_0953_9961_0362;

        #200;
        key = 128'hc07e_3a69_525b_9926_44cc_69ff_5a79_115e;
        state = 128'h0da7_180b_77fe_a2ce_630b_e06d_1831_f9a5;

        #200;
        key = 128'h0024_97ce_cce4_49d5_6309_f5b5_e487_ba6e;
        state = 128'h2ec3_51c9_db05_935d_128d_7727_c646_1d58;

        #200;
        key = 128'heff2_78e8_cfc6_4b35_864c_98c7_b1bc_b695;
        state = 128'h0e57_486f_d767_b109_b061_320e_506f_43d3;

        #200;
        key = 128'he1b6_2d11_da97_e411_f6a1_570d_7fdf_957b;
        state = 128'h5ef0_edd2_90d6_d2a9_b791_89d5_d68b_fe07;

        #200;
        key = 128'h4fb1_33b3_1703_a2e9_ca76_5647_13e9_f008;
        state = 128'hd210_1e1d_5108_d3b3_07f7_01ca_4c59_fe75;

        #200;
        key = 128'hc4e7_19f6_6fb8_90b8_2b24_8f9c_eca6_de9f;
        state = 128'h28d7_c681_bf09_dcd9_235a_f8f5_c311_5085;

        #200;
        key = 128'h6c72_510c_f42d_bae1_f25b_742a_375f_639c;
        state = 128'h4b55_1f5f_c1ec_8469_8603_6af1_73c7_6788;

        #200;
        key = 128'h4360_8a7f_4a9e_71bc_8b4e_8afd_dc1d_b2a2;
        state = 128'h7c0d_27e3_085d_424d_4a1a_be1f_7edc_ce19;

        #200;
        key = 128'h0a8c_0930_aee5_aac3_921b_d44f_971c_faa3;
        state = 128'h830d_8474_db26_e8b9_bd9e_c234_3a4f_88eb;

        #200;
        key = 128'hff02_38fa_6a73_c70e_92c6_552c_1fd7_1033;
        state = 128'h8469_b9dc_4ba3_052c_f9eb_3526_8e17_fe6b;

        #200;
        key = 128'h2a3d_3ba1_a4a1_492a_4926_0614_2253_d59e;
        state = 128'h43e6_0c33_a6d4_5055_2b73_315e_0398_7031;

        #200;
        key = 128'h0dd8_c7be_f667_800a_b07c_f18c_1691_5f2c;
        state = 128'h7e7d_ce62_261b_dd9f_44b4_3771_9f35_7f3d;

        #200;
        key = 128'hf725_01d4_0ee4_ec5c_8501_8292_4b78_98ed;
        state = 128'h394d_934e_7568_d861_0d07_a88c_6bdb_e047;

        #200;
        key = 128'h9622_daef_a4c6_14c1_7136_689d_4e8e_c75b;
        state = 128'h27dc_8188_6aa0_8672_6af0_d73b_1560_9f45;

        #200;
        key = 128'h9a3e_be48_a198_9fd1_b538_2204_fa16_b70f;
        state = 128'h763c_eb92_448b_b4cb_8887_ed46_05fb_2598;

        #200;
        key = 128'haf4c_4a6c_7794_1431_8ce4_0227_3bf8_abb0;
        state = 128'h0f5c_727c_052e_1771_cf49_cae2_cea3_c6d5;

        #200;
        key = 128'hc6a8_fdf8_23ed_2d6b_d0fd_25ef_d599_27b5;
        state = 128'h8db1_2829_7edc_2a52_c067_bbac_5352_044d;

        #200;
        key = 128'h8e82_10ff_6d7b_84b6_94f4_c29b_b18f_0363;
        state = 128'h1dc7_32ae_e293_b87d_a49b_6f0a_2010_9d41;

        #200;
        key = 128'h0c33_8a4a_c728_91da_7178_eda2_d477_b96c;
        state = 128'h9fa9_4a6b_3b96_d0c9_7d2c_e997_b7c8_15f2;

        #200;
        key = 128'h3dc5_b1e4_a4d4_c02b_d01d_3ccd_a256_95ab;
        state = 128'h3e92_a9c2_1ce3_918c_06fe_ebd5_003c_db84;

        #200;
        key = 128'hcc7a_0c0d_2bc4_c544_eef5_41c1_2b85_a9d2;
        state = 128'h1e4a_6407_3b73_9d18_434f_e386_add4_dbf6;

        #200;
        key = 128'h2a8e_5f6f_7238_94e8_d0aa_3ea1_c5c1_a221;
        state = 128'h4563_984f_5a04_62e2_9499_a454_4850_caca;

        #200;
        key = 128'h2b1a_d964_3ff2_c27d_cdf7_0e39_5405_cf22;
        state = 128'h0c68_27cc_9249_d2b4_4806_fadc_ddd9_5fb0;

        #200;
        key = 128'hf6dd_c766_9269_ad37_4375_d69f_1c09_fd97;
        state = 128'h7526_32c8_db4a_7d8f_d0fd_7e49_769b_0f31;

        #200;
        key = 128'h5766_702e_c281_58ba_67ac_820d_27f9_5e55;
        state = 128'h268c_5438_a12b_1d94_e965_cc6a_e8e8_a3f5;

        #200;
        key = 128'h53f3_abf2_7a1a_6e56_a482_1a3e_0fb3_a66f;
        state = 128'h0b9d_3780_e1e8_44ae_a01e_8e47_b1f9_b822;

        #200;
        key = 128'hab54_ed5a_21c3_2267_1245_e13a_a1aa_955f;
        state = 128'hff26_f726_bf61_9259_1c33_9264_d6af_78f2;

        #200;
        key = 128'haf24_3bcd_cdb0_e617_bdfe_a46f_5fa6_dab1;
        state = 128'h9885_2581_15c1_4794_d5ab_7ba8_f08c_6907;

        #200;
        key = 128'hc775_e37a_5b58_fada_cb8c_7b81_f03c_aa03;
        state = 128'h0118_a753_6f9f_ff21_be8e_7bee_f9c8_2e65;

        #200;
        key = 128'hf9d3_bb0f_c435_1af1_1a25_b577_ef6b_56b3;
        state = 128'h7c4d_cc2d_2c58_d645_5061_e508_c89a_3631;

        #200;
        key = 128'h14c5_7714_67e9_8e88_9987_c984_ba28_812e;
        state = 128'h0932_7a87_6bbf_f7e7_256e_7866_f8c5_d515;

        #200;
        key = 128'h127d_ca2e_6bf2_e512_3f33_c229_dda1_9b1d;
        state = 128'hbc01_266c_a318_7436_3af1_e333_d796_3daa;

        #200;
        key = 128'he696_a4b1_a534_8b0c_521d_8d55_80a5_f69a;
        state = 128'h6247_f376_d6da_f693_6ab6_05d4_f9b9_62e5;

        #200;
        key = 128'h1d56_b69d_7d2d_acd1_3aa4_3dad_46cd_1fe6;
        state = 128'h0633_2321_cd8d_1cfb_bfa7_8274_1155_e1bd;

        #200;
        key = 128'h66a2_beeb_0026_7cf2_6a7a_9b9e_c085_897c;
        state = 128'hb82c_6873_4a18_84fc_bc66_4a6c_3f2a_cb8f;

        #200;
        key = 128'h2b01_2e8f_fe6a_e767_1412_a1be_df04_b34a;
        state = 128'h0632_5671_790f_6f69_3039_697c_2302_ff35;

        #200;
        key = 128'he4c5_f551_8df4_378c_2a77_e929_c2c2_55d4;
        state = 128'h7400_a603_dde4_4aaa_975f_7730_6682_8165;

        #200;
        key = 128'hac75_cfdb_4623_b273_169f_0922_8bc1_2953;
        state = 128'h8133_bf56_c50c_4919_ea1e_94f3_c44d_7cb2;

        #200;
        key = 128'h93fa_4175_118e_b639_2199_02fa_ee84_f5ea;
        state = 128'h3a62_5ea6_aa3c_f59b_dfa3_3ee4_6add_d991;

        #200;
        key = 128'h168a_b16e_d311_b539_cb86_50f8_320d_861c;
        state = 128'h46c7_787c_e67e_07e4_60b7_5a19_de30_8c64;

        #200;
        key = 128'h7dd1_5ba8_68a6_a682_421e_a7aa_e94c_f708;
        state = 128'h2706_7ae4_c020_85aa_e1b3_ff91_14df_45ad;

        #200;
        key = 128'hef65_bb4d_8e63_ac7a_1ae9_64de_3550_02c7;
        state = 128'h7f08_c931_273b_7e32_dc69_f30a_485c_53cf;

        #200;
        key = 128'h01b5_8022_801b_477d_5bff_38eb_433d_c67b;
        state = 128'hd50a_90a9_3306_9842_41fe_9238_07d6_4a01;

        #200;
        key = 128'h904b_62bf_8b73_d9f2_9d13_6f03_c7ab_ea3d;
        state = 128'h1a96_a8d7_d4e9_b265_4b4e_63fc_1896_ff16;

        #200;
        key = 128'hb861_2d9e_c952_5e17_0c92_578d_f31a_2e08;
        state = 128'h72ba_8a53_72c5_a65e_8d86_cbdc_6e12_511f;

        #200;
        key = 128'h66b1_7d40_9754_3b55_6bff_1d5e_58bf_faf6;
        state = 128'he15b_f2fb_f9e0_789b_4302_9057_9091_a1ce;

        #200;
        key = 128'hd86a_25d4_d2f1_73fe_99dd_92d4_9f58_0dad;
        state = 128'h1327_3d1b_7b8b_f953_6e1f_ef34_8272_3ef4;

        #200;
        key = 128'h31c4_1bc4_f1cb_92d8_41ca_9b33_5f83_78bf;
        state = 128'h496b_490f_7ef5_8fe3_1ea9_f9f0_cd2e_b600;

        #200;
        key = 128'h14bf_1625_c091_feef_576e_9233_6823_b5bf;
        state = 128'he53a_213f_1107_0003_1efa_1462_8042_efc7;

        #200;
        key = 128'h7abb_ab12_9fb2_5880_f512_95b2_8b77_6116;
        state = 128'h1f2c_fea4_24cd_5239_8ac3_02d5_e463_d173;

        #200;
        key = 128'hbfc3_e09e_34c9_9498_70f1_aeee_4e5a_5598;
        state = 128'hce7b_cf12_2a5e_2d70_727b_3632_0c84_f766;

        #200;
        key = 128'hcb84_8189_7fa7_4f95_6174_53ab_e1e2_8958;
        state = 128'h49b2_2de2_639a_6f5d_5b95_bb0e_68e0_2383;

        #200;
        key = 128'ha0ff_f91d_746c_f3e2_f3f7_958f_e77f_6c78;
        state = 128'he505_6037_cdfe_e0e2_c242_0568_c6a5_f834;

        #200;
        key = 128'h125a_9729_9c8e_45b2_3a02_544a_425b_b2f2;
        state = 128'ha053_2ae4_eb05_1d3c_4d8a_e2f1_a37e_9ef7;

        #200;
        key = 128'ha088_d577_222c_292e_b928_55e5_5c89_6b8f;
        state = 128'h148e_2ed1_eefb_b390_175a_3cef_fccd_9458;

        #200;
        key = 128'hdffe_c22a_d4b3_07aa_abe7_ea3c_716c_6196;
        state = 128'h0e0d_3a7b_e3b2_5341_045a_705a_8dbe_ebf5;

        #200;
        key = 128'hd45d_db4c_cfbb_94fb_9759_9ea0_61f3_1d9c;
        state = 128'he61e_aafa_858f_f293_ec48_8c74_d4b0_b7b3;

        #200;
        key = 128'h1550_449f_1cbc_98e7_35e5_7ca4_cbb8_83bd;
        state = 128'h20e5_db93_7cbd_9f94_02c7_425f_0c60_4122;

        #200;
        key = 128'hbcb5_0754_4b9f_1c4a_8d35_37cb_1f47_62b0;
        state = 128'h95e6_27b4_f7ba_754f_dbe3_7960_87b9_4688;

        #200;
        key = 128'h370a_3e69_f814_4ba4_240a_1c51_4bdb_ec62;
        state = 128'h5fe4_9d6f_7a32_af83_3f19_2742_71ac_53fd;

        #200;
        key = 128'hbdd1_435d_a21c_58f0_ca5d_afbe_00a9_b407;
        state = 128'h13ca_4afb_2264_957c_a802_0ed8_b52e_86f6;

        #200;
        key = 128'h92b4_b175_6a2d_068a_0539_6f9d_c49c_cf0c;
        state = 128'h03ad_9d07_6e6e_3c1f_e01e_e764_b439_9525;

        #200;
        key = 128'h16dc_04fd_606d_990d_ed3d_4810_dfc6_96e9;
        state = 128'h58df_5cc7_56a5_8a0d_5fd8_19aa_ebb7_679c;

        #200;
        key = 128'h55b3_0dd0_d267_4ed6_cb77_8785_3843_ccdc;
        state = 128'h7788_29c9_4fee_bec1_76e7_5d8c_6603_c508;

        #200;
        key = 128'h206d_3285_2b73_574e_c039_a552_49c9_3ada;
        state = 128'he1e9_9c15_1747_b763_ed66_bb47_17fe_a84f;

        #200;
        key = 128'h8e24_2c85_1712_646f_efb7_ddc5_30d8_dec9;
        state = 128'hb499_773a_787e_fe4c_1e32_c218_7c49_6a6e;

        #200;
        key = 128'hddec_9e77_2880_3eb8_7f8e_9156_4e64_315f;
        state = 128'h7662_df4c_b296_162d_d186_b869_a95c_b0cc;

        #200;
        key = 128'hcb64_1b64_19ef_1cab_4cbb_27f9_fa15_9f45;
        state = 128'heef5_335e_e0a9_85b5_3c51_056a_4175_c71f;

        #200;
        key = 128'hda75_75a4_d2f6_3133_d4ea_6e46_1dac_7e20;
        state = 128'hef97_f4d9_9683_06ef_552c_8154_7f62_5cd0;

        #200;
        key = 128'h5c30_13d0_9cdc_1e7f_9bf8_aa1f_c2aa_d7e6;
        state = 128'hda6c_f173_b11e_b24d_2663_1717_5dc1_5334;

        #200;
        key = 128'hdb17_529a_b45b_8919_b26e_4047_a7ca_9edb;
        state = 128'ha1c7_d7d4_3a4d_7431_0795_8a51_3dd0_1d52;

        #200;
        key = 128'ha6c1_609e_4bef_3222_2d37_93cf_200c_ce1b;
        state = 128'hd8ca_03fc_f557_bf2e_8720_9473_d6f6_ddfd;

        #200;
        key = 128'h7916_c410_a264_8aca_b57a_f0e2_2253_7e46;
        state = 128'hba25_f596_8b01_99d9_cb23_4e74_4696_b3ea;

        #200;
        key = 128'hfc05_57fe_9a59_bb66_8aff_c83a_6564_27a3;
        state = 128'h69a9_ee1f_04cf_b471_8f50_8244_714a_bde8;

        #200;
        key = 128'h3a3a_6add_bca2_e8cd_77c4_cdd3_a47c_f87f;
        state = 128'h4d98_2438_bd88_19f4_9d7f_7f79_3739_0a20;

        #200;
        key = 128'h1389_afb5_0ed9_18ca_3cf9_dbc9_a0b8_5669;
        state = 128'hedbd_da29_9e87_1e98_3d19_6b68_86a7_058b;

        #200;
        key = 128'h6e70_7f5f_1b68_957e_1210_e25d_a009_ef81;
        state = 128'h5f08_a9ed_ad66_0826_0ad4_ec57_e71d_fc10;

        #200;
        key = 128'hd3e3_2421_dba5_6eda_a903_c32e_63b5_d222;
        state = 128'h0781_b04d_4b89_3d19_3315_e82b_a90d_9cdf;

        #200;
        key = 128'hd1bc_59f5_2fed_7bd4_19d1_2ef8_3614_da0f;
        state = 128'h8ccf_b42c_ee18_46ab_01be_bf50_60cf_adaa;

        #200;
        key = 128'h3788_ef14_f267_b791_fc2a_cf86_6a40_2510;
        state = 128'hcdcf_457f_c04b_a058_8f26_32c6_34fd_b91e;

        #200;
        key = 128'h8496_b23f_6901_343c_2257_7806_817c_87b9;
        state = 128'hb695_ac88_f17e_80c2_8d81_775e_8d96_5510;

        #200;
        key = 128'h395b_cc7d_9fcf_e86a_8a20_8099_558f_8340;
        state = 128'h5caa_7e93_6b31_4e46_a728_98c9_b1e5_e21b;

        #200;
        key = 128'hf3aa_b9a5_762b_af8c_f8b9_c809_8b6f_3690;
        state = 128'h0bd1_e040_6304_578c_f077_0fb3_1772_41ef;

        #200;
        key = 128'h4f1d_a2d7_6d68_7f2b_e7a1_dd56_eba5_2cdc;
        state = 128'haa32_ba32_e023_68a8_45b0_8102_5579_32a9;

        #200;
        key = 128'hfa04_378b_a9c3_5501_621e_8c0a_4334_3e3e;
        state = 128'hc1c1_a533_f3f8_7dce_b335_aca3_44bd_2ca2;

        #200;
        key = 128'h8dcd_54ac_b19a_c12b_7ddc_04d4_dfe4_4c07;
        state = 128'h005b_0452_ccdb_13e0_e5ab_8606_944c_7edc;

        #200;
        key = 128'h3cac_5746_2c7b_6912_8075_f000_a417_335a;
        state = 128'h0d9e_91cb_1f5e_99ea_e09e_7f83_93ce_7745;

        #200;
        key = 128'h7698_f8ed_61bc_9702_daf1_4e3c_84dd_511e;
        state = 128'h58b2_fdfc_626a_fc3b_5b0e_7bd2_ee03_09ba;

        #200;
        key = 128'h93ab_79bb_d059_a78e_188d_3c12_3c3d_8522;
        state = 128'h73d3_ebb3_5eaf_6b3a_22fd_f3f5_5017_db4e;

        #200;
        key = 128'h96d6_ef07_d8b6_e2ce_1274_9a38_4d14_1020;
        state = 128'h8bdd_b352_9d24_8983_f891_5cb5_c974_240c;

        #200;
        key = 128'h14be_011b_08b8_144c_772e_2736_db33_351d;
        state = 128'h7d9c_697d_54fe_0462_f8ff_4836_c60f_8c0d;

        #200;
        key = 128'h8dfd_22d5_e23f_2afc_692a_20c6_93c5_d4e1;
        state = 128'hdede_6820_ff44_9d5f_62ce_a2c1_4e4b_ab86;

        #200;
        key = 128'h277f_8904_8c8d_e80e_39d6_fa7b_9eb3_2ef8;
        state = 128'h6187_292b_ef8e_3115_ab5a_d126_91fb_fbd2;

        #200;
        key = 128'h2c72_92c3_f719_8c28_dbdd_2c80_0b56_b1be;
        state = 128'hfc27_4b76_5d44_a121_06cc_59c9_2ff0_d3f0;

        #200;
        key = 128'hf6a2_4787_6811_cd52_db92_868a_491e_1840;
        state = 128'h47f0_464c_031e_00ea_a779_76a3_e741_d7a8;

        #200;
        key = 128'hbf92_42f1_8964_96d2_4495_bb9d_d2d7_23d8;
        state = 128'h1f32_2764_27c3_8cab_99d3_d21a_beaf_7f72;

        #200;
        key = 128'h3ed4_e12c_24da_f775_b855_0e4e_81ad_9634;
        state = 128'hd731_bbde_205a_8695_5348_f96f_250a_ecda;

        #200;
        key = 128'ha1bf_3519_305b_4a07_c2bc_4dda_cd97_6078;
        state = 128'hd205_c4a1_f343_dae5_4ec0_a015_129a_5b53;

        #200;
        key = 128'hbe2f_562b_7356_7e5e_0da9_30c5_6f99_c35f;
        state = 128'h4a6a_780c_68e0_7c66_6485_1b35_ec88_c7b2;

        #200;
        key = 128'hbe2a_e708_ea13_9d57_c764_a6ac_0031_1dc9;
        state = 128'h943f_fe65_2ce0_c052_8522_54d8_5178_32e2;

        #200;
        key = 128'he04e_b7b2_a35f_06cd_fd8d_0f2d_dd91_aef8;
        state = 128'h8504_6fca_40aa_fa02_370e_aa43_361c_1707;

        #200;
        key = 128'h8122_a195_47ce_6738_37a4_efa7_2f0a_caf8;
        state = 128'haec7_7bf4_a743_32ab_d7ed_df63_22e8_5a47;

        #200;
        key = 128'ha760_1530_d3c2_64ba_4ca4_1e8b_037f_7b46;
        state = 128'h48bd_c944_eab8_37af_66f4_3877_4689_f3cb;

        #200;
        key = 128'h92b8_ac86_638d_2546_ae1a_e248_ffcf_4740;
        state = 128'h5d31_9b15_ec99_bebe_1bad_0e58_736f_cc36;

        #200;
        key = 128'h72e3_745c_ae90_06cb_1b98_9063_4b04_9953;
        state = 128'h1458_f89f_a1c5_3faa_5eac_a584_2449_02d0;

        #200;
        key = 128'h33d4_9334_936a_dd9d_fe68_caa8_d0ac_e7e8;
        state = 128'ha166_0e00_6d66_a7ca_4af1_df63_3a27_0207;

        #200;
        key = 128'h810e_8f08_c40e_fe12_0e80_fa00_b4c1_6143;
        state = 128'h4e8c_3426_0ddb_c2af_d576_1918_e91a_603d;

        #200;
        key = 128'h7dc9_36fa_2023_7088_e6c6_e97d_1c4d_aa98;
        state = 128'h6da4_0a01_4d19_040b_2110_d328_ba9f_1d67;

        #200;
        key = 128'h69bf_960a_c18a_0d93_9f8e_64f8_88f2_b0c4;
        state = 128'hc9fa_dd09_95be_bfcd_2d6a_7178_0476_1ce7;

        #200;
        key = 128'h0546_79b7_a689_d6a5_5256_a32b_92d0_3b54;
        state = 128'h91ce_1c1d_e490_f6ba_0e46_4dc2_db2f_92b9;

        #200;
        key = 128'h4631_abd0_1509_3ec9_4b57_5038_8927_1122;
        state = 128'haf14_4b47_93d0_d7a0_a9b0_7e85_58df_9f20;

        #200;
        key = 128'hce7f_bf13_2fa8_dd66_2819_ab66_6431_7449;
        state = 128'h888a_d3eb_ba16_12c1_9605_6ea0_373e_7018;

        #200;
        key = 128'h3b98_9ab4_c898_47f0_8d7a_3ce6_02de_b6d7;
        state = 128'ha9e3_81a2_f107_9af1_7732_a1ae_b9b5_d001;

        #200;
        key = 128'h55ec_8e61_1b02_3404_cb4d_cde3_5fbc_82f4;
        state = 128'h6092_a134_523a_63cd_6b2a_a349_339e_7d43;

        #200;
        key = 128'heca8_aa1e_64a0_d6cf_7af4_a117_8cad_fc5f;
        state = 128'h4657_801c_3bcf_19b7_2e22_d9ba_b827_6f27;

        #200;
        key = 128'h82ad_c793_9dc2_00b7_792a_8595_c8b8_4895;
        state = 128'h1771_d108_3924_3876_d414_442b_e4e0_0bd0;

        #200;
        key = 128'h845a_ce87_e64a_cd0e_ca73_c4a5_c446_9e0e;
        state = 128'he079_db11_5b46_9e95_163b_acf7_98da_c3fb;

        #200;
        key = 128'h91d7_4797_f9ab_2a84_d75d_3c58_ed25_26ce;
        state = 128'hecd1_3654_34aa_f305_15cf_9484_2211_b550;

        #200;
        key = 128'h20d8_e62f_74a7_9746_f0da_c2e1_2ca2_136f;
        state = 128'h9ecd_d399_352e_cb38_0f16_699a_bc46_e105;

        #200;
        key = 128'hde93_59ba_de1a_2303_7e28_60c7_f701_d607;
        state = 128'hb880_9c19_a936_fce0_aed2_8faa_3bf6_eae3;

        #200;
        key = 128'h8cb5_7cae_233a_5f17_ef52_bea3_b448_2272;
        state = 128'h883f_665e_f222_f9ad_892a_8a77_79a1_aa09;

        #200;
        key = 128'hea71_2b13_56d4_fc77_3f1b_9e36_22c1_9dd9;
        state = 128'h743e_8aa9_54b4_3e41_8f3c_572a_a9f5_753b;

        #200;
        key = 128'h213e_bccb_6471_5134_648e_1d35_705d_5fb8;
        state = 128'hef7b_993a_e202_dea0_16fe_b30a_2960_cb28;

        #200;
        key = 128'he2b6_d415_0921_6c68_b504_562f_4cbf_e001;
        state = 128'hcfd4_36e1_68d0_a370_cf3c_46d9_1300_2a52;

        #200;
        key = 128'he45d_52f3_7a63_cfad_ae14_df3b_bcd1_77ea;
        state = 128'h80de_5512_aa19_c762_9b44_e274_35ce_8c74;

        #200;
        key = 128'hcf44_49fe_f135_e3af_6fcd_3857_add7_0303;
        state = 128'hd75b_b558_997f_4d85_b81a_24c8_ab58_7349;

        #200;
        key = 128'h8eeb_79f6_1af3_74d6_a0cb_4bf4_17f6_36f8;
        state = 128'hcd85_a091_97cd_2713_2a8c_a4f0_af07_56c2;

        #200;
        key = 128'h9fbf_3df1_e2a0_2674_f95e_1b9c_733a_138d;
        state = 128'h705a_bd1c_cc3f_a28f_d815_cf49_e4fa_a7f5;

        #200;
        key = 128'h7255_105b_5e61_76ab_655a_745d_f7dc_dc81;
        state = 128'h8bb6_7540_bd6e_b382_102d_2dc2_6ca6_8b56;

        #200;
        key = 128'ha149_3694_e2d0_27be_7dec_13d0_5362_cc59;
        state = 128'h1cfb_bd4b_771b_52b7_0f7a_b087_da6a_7fa0;

        #200;
        key = 128'hfa6b_f28e_e136_9a6f_63e9_f6af_7b99_f354;
        state = 128'hf996_a8d1_efec_e742_09ec_2af6_f79a_ebf2;

        #200;
        key = 128'hea7a_4eeb_6b9b_7a14_5894_6caf_d70d_2e8d;
        state = 128'h4262_f948_eae6_ae0a_a8b6_2607_f8c6_5d39;

        #200;
        key = 128'h17c8_3b19_c262_0e28_9db9_99d1_9041_678e;
        state = 128'h144c_c1db_09e7_20b7_4d1c_af5d_ce55_d492;

        #200;
        key = 128'h66e3_9842_6e86_cdf7_ad1b_6e65_d35b_cadc;
        state = 128'h98d0_af06_59d3_19d3_55bc_6680_ec4e_48a5;

        #200;
        key = 128'h2907_abb4_2053_3e9f_dcbe_a4a7_d4e0_716c;
        state = 128'h3db9_d024_9be3_2d84_7197_8bff_6721_b993;

        #200;
        key = 128'he577_428a_d7dc_5d20_4a5b_edc4_bb7d_a44b;
        state = 128'h9ef3_73ec_501b_2a28_f09c_e281_c675_1440;

        #200;
        key = 128'h7c75_5851_1d2c_6a2d_20a8_7a4e_605f_3601;
        state = 128'h2768_6be2_149a_16bc_f6a5_52e7_f8d0_b931;

        #200;
        key = 128'hef45_3bcc_b0b8_42bd_f848_068e_b329_ab8e;
        state = 128'h4fd0_39db_73f1_9a6d_2ffd_7e09_b75e_4a33;

        #200;
        key = 128'hdf6a_66b2_a501_badf_7169_eb79_8eb7_9e93;
        state = 128'he7d8_757f_9b45_ebb1_321a_dc5c_47ea_aa0d;

        #200;
        key = 128'h3e8f_2781_68d2_7a14_6812_bd74_2617_109d;
        state = 128'hd873_8e09_b8d6_51c9_9d0f_8314_c087_e3be;

        #200;
        key = 128'h1051_1b57_e142_715f_5d4f_56cd_4db7_c29e;
        state = 128'h602a_133e_4df9_b4a5_e5bd_40ea_fa45_ecda;

        #200;
        key = 128'h7147_2acb_91ff_798b_8d46_92fe_23c1_bee5;
        state = 128'h71c0_c9ce_2e19_acf3_f14e_6272_f78d_778c;

        #200;
        key = 128'ha144_2243_2e59_3be4_8ceb_2ff6_6daf_cd4a;
        state = 128'ha758_fd07_12e4_8bd4_d2d7_fbc8_192b_a63a;

        #200;
        key = 128'h96f1_c4b8_dac2_fd5f_5e16_5c52_3380_59d6;
        state = 128'h53f8_ffd4_51f2_ebca_ec31_afab_a8ef_b6da;

        #200;
        key = 128'hcb13_67c8_1f48_237f_a0fc_3c9e_b15d_85d3;
        state = 128'hb93a_8401_763f_079c_b3b5_4ee9_271f_9d00;

        #200;
        key = 128'h1d95_e3c4_5e62_dd9a_143e_ec95_e9c8_0971;
        state = 128'hc855_ff97_ba04_60fa_07b5_6c4f_864e_c665;

        #200;
        key = 128'h819a_eb69_1afb_b06c_eee5_c291_34e8_dcdc;
        state = 128'he366_4ae5_aafb_4e4c_7d60_e41c_67e9_12ce;

        #200;
        key = 128'h00ea_6ba2_a0a7_4a7e_9aa8_ed2a_343e_3a29;
        state = 128'h51bd_11b6_9caa_69ec_e028_4ea9_5d17_0627;

        #200;
        key = 128'hcb92_b401_8a4b_c72a_bc11_0995_74b4_01c2;
        state = 128'hf575_4cf0_ccd5_7fe7_39d9_ccce_4016_92d8;

        #200;
        key = 128'headb_09bb_f306_a7ac_ab4f_900c_5d25_a52e;
        state = 128'h2e77_17ad_126e_d3ce_0228_32a0_0a10_17f1;

        #200;
        key = 128'h5eec_02d5_3ae2_19a5_848a_afba_6aa5_2693;
        state = 128'h4e61_9740_5aef_cfb6_8423_2870_c9f5_3a44;

        #200;
        key = 128'h5ab6_525f_39a7_c9ca_1184_7ad0_3231_d430;
        state = 128'h6703_9d82_f93c_735c_8354_9e39_1fa2_f81c;

        #200;
        key = 128'h35b7_2375_d670_21cf_ec5a_7814_9b7f_0c66;
        state = 128'hfcca_bfe1_8640_9a83_470c_69a3_1679_3d75;

        #200;
        key = 128'h1887_05da_824f_39ec_542f_a05c_b0ef_ce90;
        state = 128'h8222_7679_2184_5c5a_9b11_e273_b81a_c88a;

        #200;
        key = 128'h81d9_4314_494f_dc8b_d028_2d3a_2531_512e;
        state = 128'h8543_64dd_afda_b0b3_32fc_5543_87fa_c0af;

        #200;
        key = 128'h97ca_adab_b0ea_0bdd_f238_c6ef_2c07_e6fb;
        state = 128'h6144_92e3_cd48_2c87_a007_3b8d_37a8_a0f1;

        #200;
        key = 128'h3237_748e_dbf9_278e_ead9_cddb_8de1_7608;
        state = 128'hf97a_2ff3_d03b_b50f_b2ce_f008_81a0_08ef;

        #200;
        key = 128'h587e_76ea_de31_c92e_0264_bca9_eb94_2c13;
        state = 128'h9216_1a3c_8a7f_a2bc_8889_6f0c_63f3_928b;

        #200;
        key = 128'hc194_3291_b25d_54d0_faf0_d972_791b_2d43;
        state = 128'hafbf_2a02_a346_73f4_5033_0d57_034a_1fde;

        #200;
        key = 128'h9890_4d8e_646f_811c_8568_343e_722c_3c3a;
        state = 128'hbf2c_e9f6_08d7_15bf_2235_fb51_2b70_8921;

        #200;
        key = 128'hd94f_11f2_29f5_a433_e7a6_c5e2_439a_2b1c;
        state = 128'hdf13_0d8e_7047_5306_bd4b_4d57_1dba_8743;

        #200;
        key = 128'h9e28_a19d_b775_e035_dce7_d5e8_8782_e03f;
        state = 128'h30c6_e239_6844_c5a2_190d_26e8_1272_4850;

        #200;
        key = 128'h5644_04f4_6eb1_36c3_b71e_4ea9_97cd_683b;
        state = 128'h4665_c9a8_8c9a_702f_26f0_516f_6069_b718;

        #200;
        key = 128'h41f3_a82d_5a98_364a_eb06_f005_6686_34c6;
        state = 128'h61aa_af56_8479_d9a5_9eff_c143_0fbf_9f1f;

        #200;
        key = 128'h3828_f354_e53d_8187_f638_9313_e8b3_7e82;
        state = 128'hc27f_0260_9430_a8de_0e88_47f2_af00_9dff;

        #200;
        key = 128'h26a4_f74a_4ba7_ca27_494e_a214_927a_e355;
        state = 128'hc595_fc31_ff58_5297_3dc6_de69_199e_5e39;

        #200;
        key = 128'hf366_47cb_996a_c04c_cf8c_4d24_bd10_ed10;
        state = 128'h744e_cb2b_efa7_6166_a0ec_231d_3eb7_a2fc;

        #200;
        key = 128'h7ab1_d9b0_ab6d_978c_8f87_ebc4_a6ce_1a6d;
        state = 128'h8ec1_cb46_985a_6375_20e1_00e8_f477_8e76;

        #200;
        key = 128'h35fb_380e_c1db_0989_ebac_55f9_6363_9023;
        state = 128'h040b_5603_efc4_9973_353f_66c6_f183_786c;

        #200;
        key = 128'h60af_c746_1210_47de_e284_7e0a_afde_16bf;
        state = 128'h3007_148a_6557_deca_6ee0_950a_a329_5a94;

        #200;
        key = 128'h3c4e_ee9b_78aa_7e0b_ace3_ca1c_ce74_8d96;
        state = 128'hc8fb_bcac_0d1e_4572_ef37_6328_6e57_6d78;

        #200;
        key = 128'ha9eb_f7b1_3d78_224a_7a18_48a1_f6ca_c81b;
        state = 128'h477b_a42d_0c0d_a8e5_6d6b_61eb_7e9d_6bae;

        #200;
        key = 128'h20dc_72de_a9cb_f534_b219_93b9_b5f4_77f5;
        state = 128'hf1e6_85ea_f510_c54a_b1fc_da91_d993_72f8;

        #200;
        key = 128'h3941_d68e_0607_7403_2289_9080_407d_3420;
        state = 128'h1ec7_b44e_e283_1c96_566f_c43f_e5c7_cac5;

        #200;
        key = 128'h1fe4_9eaf_ec8b_b197_fdfb_37dd_496c_b319;
        state = 128'hcaef_6139_68ac_eba1_d469_2ffe_2a84_59fe;

        #200;
        key = 128'h5843_1b46_bf1e_8fc2_7714_7069_c38d_d4b5;
        state = 128'h0f7d_37ea_b6b6_6829_c880_c5e3_cb9f_a25f;

        #200;
        key = 128'hed59_408c_c83d_ca8a_6142_133c_70e4_6b51;
        state = 128'hcfa3_427c_98b6_f76c_99b4_1e8a_59c9_52d6;

        #200;
        key = 128'h0e78_1e66_c913_9ec4_5aae_fb8f_b575_d0b5;
        state = 128'h0b6d_2eab_eddb_91b1_14b7_07d6_64a1_72d1;

        #200;
        key = 128'h7050_63f8_49d1_7cd2_77d9_53e3_d432_895b;
        state = 128'h8068_dd23_09c0_ae4b_534f_36b7_e917_bef7;

        #200;
        key = 128'h17ad_bd50_f385_c653_0a53_ec5f_0805_1c5f;
        state = 128'h97e5_172f_6850_dc37_ee4f_5879_dc1e_87c4;

        #200;
        key = 128'h5dab_82d7_fec9_cac0_dc69_cf6c_e3ce_d86e;
        state = 128'hbb9b_91d7_81f7_c737_1f5f_4f0f_2893_0233;

        #200;
        key = 128'h464a_eaab_7c23_35a4_a5f4_bc15_1c82_d07a;
        state = 128'h7fa5_488c_6f4b_8028_6814_dbd1_57c0_58e0;

        #200;
        key = 128'h31ec_1461_c2ef_87d4_346f_3796_b688_49c3;
        state = 128'h3081_f961_9397_8dba_2faa_3c21_c149_0aa1;

        #200;
        key = 128'hecf4_ea70_a3a5_916e_6f0a_5d0b_4b0d_ae8a;
        state = 128'hd52c_a52c_0f0c_4867_d7ca_e00b_c7b0_3d36;

        #200;
        key = 128'h0b4a_8011_b271_bcb0_2971_f368_235f_7d91;
        state = 128'ha7d8_9c0a_651a_28d9_2562_32b4_97f9_ab89;

        #200;
        key = 128'h07db_1c53_924e_5c0d_1f46_2c77_27d1_6843;
        state = 128'h392b_78c8_03c1_fcf5_b87f_95c9_b9fb_a168;

        #200;
        key = 128'hee60_8093_8c63_00d0_3f8c_747d_1c17_1c2e;
        state = 128'he276_f2a6_f904_47ab_94c8_0d4e_d444_fbb2;

        #200;
        key = 128'he5a0_6b9c_6829_bd6d_2776_dce3_a886_1ad6;
        state = 128'h1de4_9d65_6178_2390_1735_68ed_42d5_bb54;

        #200;
        key = 128'h517a_52f0_287f_4d18_aa86_af02_a415_60dc;
        state = 128'hc8e9_571b_ceee_ac05_42da_92d6_6c91_5d90;

        #200;
        key = 128'hd90f_e02f_66c9_eb40_5ae7_af48_5a19_ed75;
        state = 128'h965f_4e09_bc44_db87_82ab_44f8_f871_01ae;

        #200;
        key = 128'hd549_e5d6_af0f_b35b_22cc_cc11_cf37_d015;
        state = 128'h2020_29bb_96a7_5f2f_cf42_c7d7_ea59_3e88;

        #200;
        key = 128'h10e8_0872_1a39_aaeb_d3d5_35f3_70ec_6703;
        state = 128'hae08_7b61_527d_48a0_b933_1fc5_7587_926b;

        #200;
        key = 128'h216b_e722_52ae_a974_75b3_a570_fa58_e3a3;
        state = 128'h89f4_82d7_bda1_8d4c_e820_b5ae_2519_85d5;

        #200;
        key = 128'h6e41_8d77_cdbd_e84f_6c96_60a3_67cc_5c8b;
        state = 128'h9f6b_eb47_96e4_90ea_b5d9_abed_0e5d_6e4a;

        #200;
        key = 128'hc43a_5427_9856_632f_eca4_7ccf_462e_b24b;
        state = 128'h2229_e490_b3bc_7e28_e401_ced6_f062_ea8a;

        #200;
        key = 128'h5974_8c2e_ad27_f329_80ac_67f9_67c5_bd77;
        state = 128'hd4eb_acf2_48fb_98d5_9b22_c4ad_a2aa_d3d6;

        #200;
        key = 128'h3bdb_7e8e_8427_d018_449a_2ca3_ada5_2502;
        state = 128'he188_78b6_ca87_8338_2223_0683_feb7_d0cd;

        #200;
        key = 128'hcea5_ca9b_cc3b_41e0_1983_5884_b08e_0bea;
        state = 128'ha561_8519_bd19_1359_8c19_b0b9_e004_8948;

        #200;
        key = 128'h276a_4dac_2d37_94f6_e7e2_be5f_1b3a_08ca;
        state = 128'h42f3_0263_3ea6_e1cf_a570_d124_5f2f_217e;

        #200;
        key = 128'hcf92_d016_06a6_3a76_4241_44ef_6b61_070d;
        state = 128'hfb33_59f9_7ac4_8c88_d1fb_4360_918b_69bd;

        #200;
        key = 128'h85a1_de4b_7802_c4f1_c698_e341_0f39_8b3e;
        state = 128'ha770_e66d_e864_a099_ca30_73a3_4187_9e17;

        #200;
        key = 128'h72db_151e_eab3_6dc2_e808_7c8f_d1ec_cd2a;
        state = 128'h9e73_8e53_75b5_66fd_1844_584c_e047_e65a;

        #200;
        key = 128'h6014_955b_1a95_8a06_02e9_5810_1dcd_2e12;
        state = 128'h75b8_2139_900b_1f90_f526_59cc_ac47_4935;

        #200;
        key = 128'h3bd3_906b_580e_9d51_2b79_822c_9211_6815;
        state = 128'ha4ac_23d3_88dc_7236_38d8_1218_2534_c49e;

        #200;
        key = 128'h7359_212b_e7e2_a302_3304_1be7_6c56_a271;
        state = 128'h96f7_6fcd_1c3a_da87_4178_3214_5e5c_3869;

        #200;
        key = 128'h0739_664a_0a10_f5a9_2f77_09d9_517e_5c51;
        state = 128'h46ff_2625_e10c_507f_d0db_0f06_6114_ef89;

        #200;
        key = 128'habec_b169_3926_f91a_fd1a_4458_4f43_a4b3;
        state = 128'h9a20_c3d9_b212_3437_e5af_62a0_2fa3_404b;

        #200;
        key = 128'h9dbb_08de_1011_413f_9c90_e0e1_9a11_5159;
        state = 128'h05e3_6b0d_f9e0_0a00_ba0f_efe5_14a6_184e;

        #200;
        key = 128'hbdf4_919e_796c_3bae_5236_7318_b5aa_caef;
        state = 128'h64ba_c55d_0d0f_ccf7_aa4a_5091_f30c_0744;

        #200;
        key = 128'h17ef_f948_b1bf_0068_2469_f73a_6869_5045;
        state = 128'hd88c_3b5d_d55f_a393_2a27_9cea_af77_a157;

        #200;
        key = 128'h581b_ba9c_52c6_73f6_7af9_8f51_11eb_05ad;
        state = 128'h759b_c33f_6d20_05fd_a760_77ad_adda_62f3;

        #200;
        key = 128'hdbdc_cce6_288e_035c_4229_53f4_5164_a7f0;
        state = 128'h088f_aafc_475d_9097_decc_c6d8_167e_31ec;

        #200;
        key = 128'hbfee_c374_3a53_09fe_870c_4144_4cea_1f5f;
        state = 128'h5b6c_a239_1134_47e6_811e_294f_358e_8543;

        #200;
        key = 128'ha092_c602_69c3_4b38_ff3f_0dd4_5892_b4ba;
        state = 128'he8e3_7c9f_6823_afab_bf01_ec22_7c93_cad4;

        #200;
        key = 128'h4527_89b7_be59_8e27_58c2_b7a4_5968_fc5e;
        state = 128'hd886_5f42_d122_983e_09fc_ab02_d8fe_455a;

        #200;
        key = 128'h3680_f691_753d_9ed5_3046_1250_6ad0_e822;
        state = 128'h5d37_62e4_3a51_6dc7_534d_eb60_fed7_722e;

        #200;
        key = 128'hca74_4238_ac90_0296_e9f2_689d_68d0_b005;
        state = 128'h38a1_134c_988e_17bf_a846_b08b_a67b_57c5;

        #200;
        key = 128'hf9cb_7cb3_7423_ba0d_fac5_723c_c126_9bed;
        state = 128'hf74c_4037_1e6b_36f7_0ff8_fd1f_729d_b505;

        #200;
        key = 128'h3ea2_1db6_fcb1_1947_4e1a_b33e_d0c0_c248;
        state = 128'h5055_1245_e751_7a03_a741_bbff_9ddd_8b8e;

        #200;
        key = 128'hb594_0977_c911_c1a6_6ba5_4c73_b9a8_46e9;
        state = 128'hbcec_e495_f40c_311d_d94c_49be_52af_9ef1;

        #200;
        key = 128'hf42d_241d_7cde_9ef3_8288_053b_7705_6464;
        state = 128'h18fb_ed2b_3066_a930_4d46_f8d8_732a_a708;

        #200;
        key = 128'h860c_2f8d_fdc4_7cd5_f182_9a88_f176_9369;
        state = 128'h58cc_ef75_8698_2b74_f3f6_2e5d_0b83_ceee;

        #200;
        key = 128'h758d_b4d2_9c52_1476_3ef4_3936_9edf_835c;
        state = 128'hd663_7982_8ea5_699b_29f8_bba6_1c81_b6a9;

        #200;
        key = 128'h424b_8ba0_a6a9_4926_8e7b_db63_a028_bd6d;
        state = 128'h45c8_57bd_65e9_c60a_3b26_72fa_470f_258e;

        #200;
        key = 128'h16d8_3fbe_656d_08cc_d933_c6d9_b6c0_f4a4;
        state = 128'hfe32_50a8_7447_01ac_ac3d_481f_4804_ace1;

        #200;
        key = 128'h7794_3bda_d54c_4f45_8fac_9a02_9b53_8bfd;
        state = 128'h1e1c_7011_a8fb_cb08_9ea4_141c_71f0_4605;

        #200;
        key = 128'hcb5e_c6ec_a323_879a_bd11_c12c_3e69_8f05;
        state = 128'h1275_3f6a_a4b9_fb80_5dd9_dbce_8f88_fd02;

        #200;
        key = 128'hee21_0491_a69a_8fd0_f626_d75c_bb07_4676;
        state = 128'h80a8_bd62_cf6e_9fa9_2c78_adb6_d0ad_4655;

        #200;
        key = 128'h84b9_7a40_e959_600f_2440_a4b4_44b4_ca49;
        state = 128'h5237_0dd8_ceca_99f6_15c6_8567_4c21_f44e;

        #200;
        key = 128'h2e12_dad2_fca7_9960_2a50_a94e_cbb0_ea29;
        state = 128'hfabd_71b3_6d6e_7e05_dd51_8673_24b3_e2ae;

        #200;
        key = 128'h548d_5259_6c6c_6876_366e_c9db_302d_0c80;
        state = 128'hcb1b_c095_cb73_a37a_d1f3_959d_ae9e_9bd7;

        #200;
        key = 128'h7936_04d8_10bf_50ac_639d_d849_a2da_dc5b;
        state = 128'hf901_0a01_1fe5_4695_6b80_5e33_996a_fc31;

        #200;
        key = 128'h82f2_fe3f_3362_c367_8533_91ac_2e92_e7c5;
        state = 128'h2212_db45_8820_7df1_cac8_16a9_598a_224c;

        #200;
        key = 128'h83ad_2be9_a879_15c7_50db_8e27_f657_58ad;
        state = 128'h991e_f742_972c_a0e8_0409_5a43_c8a8_3601;

        #200;
        key = 128'h690d_cecc_f988_289a_8923_7c1f_b333_ccb6;
        state = 128'ha99e_0f59_276d_1fbc_e7a8_72aa_8027_d6f6;

        #200;
        key = 128'h7b48_9e13_bf8b_1e66_e5c7_cb31_e3a6_cc3a;
        state = 128'h6ca8_331b_215b_2153_6fc2_163b_6306_8cff;

        #200;
        key = 128'h4d90_6f0f_366e_bc2f_6fff_4dae_3dfb_0f5d;
        state = 128'h0629_2788_8509_b1f1_3b2a_2657_cc5c_5e11;

        #200;
        key = 128'h7427_b39b_6d3e_a2e7_a172_732a_5981_7788;
        state = 128'h6173_43a6_f89b_92be_1123_51db_5354_c3e2;

        #200;
        key = 128'hd077_28b4_e72e_558e_5bc2_ca70_7457_a818;
        state = 128'hb556_439b_3930_35fe_dc1e_686f_b02b_88c2;

        #200;
        key = 128'h1a1b_90e4_57e0_1fa2_3553_3a7e_e4a2_c233;
        state = 128'h7941_6ee1_3c5e_6fc0_8d22_0578_c023_888b;

        #200;
        key = 128'h01df_d99b_f87e_040b_b575_9bad_ebf7_b2a8;
        state = 128'h961c_9b4b_bc63_6535_c87f_f782_3fc9_91c3;

        #200;
        key = 128'h9605_6ce3_cce5_98ff_4194_85bb_a354_5253;
        state = 128'hb451_264c_3838_40e9_afed_111c_9deb_be0f;

        #200;
        key = 128'hc20a_6fea_03ba_1308_7896_a856_1c90_fe82;
        state = 128'hc668_82f8_6377_6d95_69d5_2991_c78a_9c49;

        #200;
        key = 128'h44c1_1e41_284b_fa44_72fb_93fa_29fd_10b8;
        state = 128'h9f47_e011_3529_773f_ab87_b29d_0866_e0cf;

        #200;
        key = 128'hc871_e5e8_d69c_b2b2_bd18_45fb_6cb6_c470;
        state = 128'hc48e_09e8_70b7_b259_d1a8_7d44_4f6d_2eea;

        #200;
        key = 128'ha71c_6d3e_f148_c396_8f56_746e_e982_8851;
        state = 128'h11cb_68a9_14b6_575c_5dd0_c0e2_3ac7_7aaf;

        #200;
        key = 128'h9d27_7518_193f_c042_2980_0d6a_3577_1c19;
        state = 128'hfb7e_19b5_76dd_eea1_0c78_0b09_f394_1ff5;

        #200;
        key = 128'h453f_5e15_8985_43ee_1f59_8e5d_dc51_a35e;
        state = 128'haa11_8f31_315f_0185_e470_cfb7_a4db_353d;

        #200;
        key = 128'h7bb9_be76_0924_f35e_2eb3_591d_2759_94a8;
        state = 128'h83f4_38a0_4e6e_c1e9_ed16_da4c_3f05_5acc;

        #200;
        key = 128'hd0a9_2bc9_da48_c571_32e5_3d7b_7c64_4e6a;
        state = 128'hd98e_51f1_8359_f332_af02_2593_e985_fa9c;

        #200;
        key = 128'h0484_dc81_b8dc_088e_d2aa_2c4a_c379_4ad4;
        state = 128'hff1a_0082_935e_4723_920c_6727_067e_896b;

        #200;
        key = 128'hfd5c_ef15_bcf3_f3e4_d866_bee5_1a34_ce4d;
        state = 128'hde6c_da75_da12_0f10_4b3a_957b_21cf_14b1;

        #200;
        key = 128'h85f3_9402_03d2_3df0_95fd_3774_a095_2b50;
        state = 128'h8296_0e6e_64cb_26d9_5f87_f905_ddb5_6d95;

        #200;
        key = 128'hf374_a3be_0527_61f4_402b_d142_3b10_fcb9;
        state = 128'hc5c0_4729_360f_87d1_9b2d_0bec_b31d_2746;

        #200;
        key = 128'h8872_c33d_0b1b_b58d_b695_445c_4ed0_e904;
        state = 128'h2f4c_0711_4b8c_4fad_d60c_21fb_d3ef_2cf9;

        #200;
        key = 128'h8433_bd51_00d4_929f_2d66_3ab4_4c70_daf8;
        state = 128'hdd95_facd_4722_7344_46c8_9de3_5874_c070;

        #200;
        key = 128'h04f6_3b17_e098_2912_b8c9_c495_267c_21da;
        state = 128'h9db3_7c16_1e0c_06f1_6ef9_3ab3_a1ad_0f2f;

        #200;
        key = 128'h74fc_ce16_650c_a5d1_7094_aad9_a8ac_2419;
        state = 128'h8107_bd8d_24f4_b177_149a_fb0f_759c_5c31;

        #200;
        key = 128'h97c3_2b51_23e5_5148_095b_8d3e_308b_66b2;
        state = 128'hf80a_53eb_dc41_a4b9_08d4_69a7_ce65_4dcd;

        #200;
        key = 128'h0cd6_efe9_995f_5a51_bc8f_3b92_ea3b_4c4f;
        state = 128'hf775_c7c1_6e6f_c026_7e79_a5db_2ba3_7e0c;

        #200;
        key = 128'h8e6a_3a5b_4dd6_810a_479a_4414_cdb7_5d86;
        state = 128'h99a4_3b33_2866_9215_2f4f_8ae3_adaa_53aa;

        #200;
        key = 128'h50c6_c1f7_82b5_5d8b_307b_f136_b531_88c6;
        state = 128'h37c2_e099_384b_2f36_75fe_b5dd_ceeb_0a60;

        #200;
        key = 128'h85f1_0cc4_e55a_8594_7b2a_b7ff_3b4a_d21b;
        state = 128'h7a97_df10_4715_1258_40c3_421f_cb37_d96b;

        #200;
        key = 128'h2c59_6fec_dec4_5cbe_0dd5_7564_b968_315b;
        state = 128'hcad2_3af7_c51f_7eb0_639d_f438_bcd5_1dcf;

        #200;
        key = 128'h720f_a3a3_696d_a64f_55a7_544e_8795_ff42;
        state = 128'hfeb9_6eab_14d6_26b8_0c2b_3ca4_396b_33b8;

        #200;
        key = 128'hcaa3_6af7_ddcf_7261_2a0e_ba01_458e_e1df;
        state = 128'h894b_3be0_3b89_48bf_b852_81b1_faab_290b;

        #200;
        key = 128'h8745_5c72_8d56_844c_b983_413e_7ee6_7e0e;
        state = 128'hde5a_7147_132e_d02e_f028_11ed_33d2_6ce7;

        #200;
        key = 128'h7176_c6ce_5a33_cd85_1608_37c9_4c58_2e8b;
        state = 128'ha8d0_e77d_41d0_e4a5_3f63_cf1f_daec_d458;

        #200;
        key = 128'hcce9_6de1_824e_dd3b_5a9b_889f_18a9_5904;
        state = 128'h1b6d_f69a_0e01_ba94_651e_70e8_f553_fa41;

        #200;
        key = 128'hec94_3a6b_c290_9a84_f162_7256_be63_c44c;
        state = 128'h20dc_288b_951c_0a69_3ec5_8a0b_dc53_72d4;

        #200;
        key = 128'hc5df_4312_4b4b_fb88_0b6a_5704_cab7_fa5f;
        state = 128'hebc2_3068_1a1c_62c3_46f8_c128_f66d_1e4b;

        #200;
        key = 128'h1c94_ca74_c0b4_6d5a_6feb_f680_328e_a5c9;
        state = 128'h38cc_b19c_e463_9841_e2b5_5eee_8327_7d63;

        #200;
        key = 128'h3302_a5d9_3e6c_76e0_0602_a2a8_ee1a_e8c3;
        state = 128'h8032_7b67_c3b9_924b_5347_6539_a644_611a;

        #200;
        key = 128'he08a_5b99_6b8e_3773_87fe_e035_bb25_4628;
        state = 128'he04f_a82f_9236_dfda_6cd7_151e_357e_6579;

        #200;
        key = 128'h45fa_183e_62fd_cf07_2b44_ce68_34ee_d378;
        state = 128'h0365_5e5e_1335_33f9_a10f_14bc_a0a7_25c9;

        #200;
        key = 128'h76b1_2236_ab0d_e277_aa89_ba3d_a098_5305;
        state = 128'h4f18_9b3f_99bd_4744_a883_750e_2499_14d0;

        #200;
        key = 128'h0a1e_b60a_3f1e_fc8d_da26_c82f_8d00_552f;
        state = 128'h7dae_0677_1f27_9bee_1d1c_6999_09ff_c137;

        #200;
        key = 128'hb15c_d50b_872f_0e8c_eb36_ad3b_e636_b76d;
        state = 128'hbfb6_0e74_2e0e_c2f2_072b_93c7_baee_c058;

        #200;
        key = 128'hbd52_30aa_c055_b1b5_8b76_96f5_14c2_13e0;
        state = 128'h0208_65e8_e407_e616_3e35_ae8b_980e_f862;

        #200;
        key = 128'h03b1_ab91_af55_d8ba_174a_052e_851c_3358;
        state = 128'h1d6d_9dcd_468a_8dc2_31c7_6d9a_94aa_d3ce;

        #200;
        key = 128'he0d4_9a85_ecc8_6396_43a2_4d2d_e599_bf33;
        state = 128'h5059_aec2_a32e_6ef0_02a4_9b35_9698_ca2c;

        #200;
        key = 128'h5f4d_60e1_ad1b_cedf_b38a_20ba_f8bb_82ff;
        state = 128'hefe4_32ed_8599_35f9_f7f3_d6c4_34bb_c285;

        #200;
        key = 128'he602_68cb_4070_68a4_3585_e28a_b32a_3f0b;
        state = 128'h4dc4_1acc_fe3e_b291_7359_3a5f_8326_648d;

        #200;
        key = 128'hc8e8_5496_145a_e89c_109d_74a9_9d7a_1c76;
        state = 128'hf8b6_4d4c_0035_a082_d5b6_888e_c54b_b93c;

        #200;
        key = 128'hef16_49d1_abf3_e7fb_9606_ed54_796a_5027;
        state = 128'h25b3_f80b_93e2_fbf2_efe9_c2d1_4c87_fb8d;

        #200;
        key = 128'hb911_1954_edcc_6077_0e47_780d_ba74_d8c6;
        state = 128'he317_9885_af28_108c_b3b4_318e_3d8a_8aad;

        #200;
        key = 128'h48cf_5756_d9c9_05f7_c674_f408_2cae_9677;
        state = 128'hf1c2_5165_1ad6_53fe_4a63_8718_5629_a09c;

        #200;
        key = 128'he6b0_2978_137f_a977_b904_34e3_efe3_b909;
        state = 128'h5ced_613f_818f_8f84_0d40_8a63_5e66_cf5b;

        #200;
        key = 128'h4c59_e85a_8b84_3825_38bc_c8f5_959b_bffd;
        state = 128'h5214_bd76_65cf_6fdc_3751_5445_91e1_2937;

        #200;
        key = 128'h0f25_b374_7ae4_d668_0a8e_aa4d_b619_7f87;
        state = 128'hfe3c_1a5e_c10c_2a2c_ac83_397f_f44d_555d;

        #200;
        key = 128'h093d_621e_2c0c_d637_554b_dad7_f1a4_c6d0;
        state = 128'h6e5a_c063_3bb9_27f0_33b8_06d4_3963_6ba2;

        #200;
        key = 128'h21cd_94f9_10c3_c479_d052_005f_9fc1_055e;
        state = 128'hce50_f35d_5012_4d86_6622_cfa3_e5cb_e69b;

        #200;
        key = 128'h8afd_1576_2735_3c2c_657e_5a9c_f65b_4571;
        state = 128'h6093_18a7_20fc_092e_5e29_7795_d6d8_78f4;

        #200;
        key = 128'heeb5_492c_f100_dbcd_049d_b9dc_5827_222a;
        state = 128'h7a0d_c485_21fe_9669_921c_af25_8779_2c63;

        #200;
        key = 128'h0fc1_7ead_4d5c_7a7f_5eda_095b_c49f_9b95;
        state = 128'h5739_de6d_84d2_1627_2d38_cc53_2a66_c104;

        #200;
        key = 128'h45bb_5e69_e9a6_93cf_576a_538b_457a_def6;
        state = 128'he4e9_dd4e_877c_4146_8598_53ec_448b_6f41;

        #200;
        key = 128'he674_8777_70f0_f93a_dfb4_ba6c_c7bd_2fc1;
        state = 128'h207d_4282_af39_ac18_ab2e_70d4_dd20_f10a;

        #200;
        key = 128'h2943_333e_5a64_dad1_caac_ee22_beb5_43b6;
        state = 128'hd750_50b3_8b85_aba7_76e9_de9d_cb25_cc5f;

        #200;
        key = 128'ha42d_8b7d_41a9_9506_298c_18ab_6ce4_245c;
        state = 128'hab18_00e9_81d5_7585_f362_2299_d9e0_19ed;

        #200;
        key = 128'h4239_19e1_b23d_92c3_1221_0f87_aac7_c7fd;
        state = 128'he269_9a07_d7da_d18b_5d55_f38d_7e14_a6a4;

        #200;
        key = 128'hea9b_2a6a_e335_c6cf_04f6_420b_2a79_cd46;
        state = 128'hbeb5_bf86_3985_228e_eb35_0ae0_5fb6_85a5;

        #200;
        key = 128'h4a51_8e7e_2101_294f_ab9e_3504_4484_c107;
        state = 128'hd3dd_dae0_61d2_4562_b8e0_c64a_ddfa_a3a8;

        #200;
        key = 128'hd7af_11c8_a6cf_bdf0_4999_2efb_c213_24aa;
        state = 128'h3006_cdbb_0b55_cfac_8786_5882_bc47_1f4e;

        #200;
        key = 128'h46ac_31c1_6760_9e46_831f_3718_b422_b785;
        state = 128'hcbea_8cb3_2fd6_7472_5196_779d_ee1a_f2a0;

        #200;
        key = 128'hebf1_59c2_1ea2_21e4_a8bf_1239_301c_7f7a;
        state = 128'he181_61b0_714d_773b_3856_3597_6d6e_f9f0;

        #200;
        key = 128'h3328_3929_b2ff_e82d_be41_01de_1d63_9f46;
        state = 128'h3ce1_9259_16fc_e8d6_ff53_0fcb_4b09_4a66;

        #200;
        key = 128'h62e3_a53a_554e_1c71_7b06_dad0_70ba_42fd;
        state = 128'h406e_0e4d_b776_09b3_8fd6_179d_6a57_514a;

        #200;
        key = 128'h584a_f828_7c5d_0f26_66eb_6502_b4a0_f529;
        state = 128'hb17c_e43c_b198_5f23_1140_b4c4_843a_5387;

        #200;
        key = 128'hfaaf_7058_8378_5dc7_756a_c487_4eae_d6cd;
        state = 128'hf6f3_f8ee_e34c_6dc8_3269_f25d_1b27_4d1c;

        #200;
        key = 128'h97c6_3fe4_db3d_3934_236b_c825_ae7d_f057;
        state = 128'h22fb_38bd_ac2a_e29b_a912_ad2a_be1e_0711;

        #200;
        key = 128'h33f6_cf0f_822f_1d53_293c_9627_f5c4_bbc7;
        state = 128'h6f1e_74b6_fba4_19aa_48c8_ecac_6546_9da6;

        #200;
        key = 128'h98b4_5ad2_44a1_1d69_56bc_b5c7_5166_79bb;
        state = 128'h1b58_9965_4dc5_d664_e25a_3ccc_35ef_431a;

        #200;
        key = 128'hc022_dfc0_00f8_f465_d6d9_59b3_eb7f_7d4a;
        state = 128'h0ec4_2a6c_55c2_768a_e8d2_d436_b787_2056;

        #200;
        key = 128'h56b5_7f2c_9ff7_61f4_d539_2e84_4383_b57c;
        state = 128'h3500_3fa9_225b_dd8c_38af_0d54_1cff_cab6;

        #200;
        key = 128'hbd24_44af_b58c_904a_8f0e_a7be_2bca_4d11;
        state = 128'h5329_2abf_2f0b_5f4d_129b_6a5d_4867_fae2;

        #200;
        key = 128'h16fd_e8f4_1169_fec7_fe1b_a8ce_db56_a743;
        state = 128'h9712_16f5_18d5_df2b_61a5_73ac_fd8c_7f16;

        #200;
        key = 128'h3cb0_ff52_d9a0_8fbb_f561_1595_67ec_2f4b;
        state = 128'h1728_5197_82b9_21a8_f47b_61b5_181a_2cb9;

        #200;
        key = 128'ha5f0_6766_8b4d_79a8_1c89_448b_f38a_3fb5;
        state = 128'h4317_fe0b_04a3_d6ec_1357_8b74_35a5_7088;

        #200;
        key = 128'h59be_1fbd_f0b4_f755_5afd_461e_0fac_f1a1;
        state = 128'h5c95_5ca1_5acf_affd_da5b_d121_a97f_936b;

        #200;
        key = 128'h4fe5_a695_ce80_bc39_f27f_e78a_93ac_0ada;
        state = 128'hff27_a0b0_04cd_8711_5dab_aa59_7a66_a4cd;

        #200;
        key = 128'h5913_371d_21ab_690f_9022_60b5_87d5_142d;
        state = 128'h4efb_19aa_4ac1_72b6_2454_2081_533a_d9f5;

        #200;
        key = 128'h59bf_8da1_99a9_5c2f_5dfa_dc5e_33f1_c01f;
        state = 128'hfcea_fa01_c2f0_0e37_ffc9_50cc_0995_f086;

        #200;
        key = 128'hbdb2_ea78_d4af_89d6_100d_b7bb_f56b_dae1;
        state = 128'he175_a4ec_c487_b00a_9fa1_679e_534e_4355;

        #200;
        key = 128'h40c2_5df2_4345_043a_1aa3_9733_fe62_fb56;
        state = 128'h385b_761b_f900_dcb5_e1cb_442e_11fe_eebf;

        #200;
        key = 128'h7841_badf_53ca_b3d1_fbef_ac56_7d80_e8b3;
        state = 128'h7f64_26a7_6f47_3872_635b_a5fc_9db2_a8b5;

        #200;
        key = 128'hcf06_7fe2_f0c7_5897_d80c_e1e5_ba89_64a9;
        state = 128'h380d_9986_f93e_1009_8a6a_e39d_3064_8895;

        #200;
        key = 128'h1bd8_3381_82ec_20d9_687e_0e4e_aa20_0f69;
        state = 128'h7d0f_3adb_ae3f_124f_0286_6227_75eb_d070;

        #200;
        key = 128'h70dc_4323_7426_a227_e11a_48f8_8355_5195;
        state = 128'h4b35_5fea_a370_1a95_9b22_9047_4c9c_a8dc;

        #200;
        key = 128'h5a1a_8320_5c3c_d182_e0c6_2287_ed68_ad72;
        state = 128'he16f_b99b_813e_7758_1e34_2f6a_66e6_e060;

        #200;
        key = 128'h4154_79e7_1518_c74b_f96e_9006_64e9_3a07;
        state = 128'h993d_5a9b_0f7a_6d2f_9e3f_50ce_4b6f_89c3;

        #200;
        key = 128'he8b9_bfd5_2596_fd56_55ac_4e51_fba9_49bb;
        state = 128'h8d21_cacc_d847_0153_786f_587f_b2fd_d478;

        #200;
        key = 128'h25d0_a752_1cf3_f5db_e462_ed1c_7809_8fca;
        state = 128'h81cd_f248_23fa_22f7_ac40_13c0_1cc8_ea94;

        #200;
        key = 128'had80_57b2_ff6b_f978_b0ee_d5ca_eb9d_72a9;
        state = 128'hc31d_7337_818b_3657_c9b9_490b_7288_4eff;

        #200;
        key = 128'h7c63_862c_b2c0_8a33_1ed1_99d2_dc61_75b5;
        state = 128'h2b4d_6386_1e12_321f_2de2_f24d_4047_e721;

        #200;
        key = 128'h76ab_be0b_2a20_97a7_a55b_ec0e_42ed_b1ba;
        state = 128'h1b0d_45b8_ae49_0728_72dc_3ca1_c689_c022;

        #200;
        key = 128'h86a9_a44b_68e9_3e97_33c7_319e_2dc2_40e2;
        state = 128'h7daa_7c5b_4cc4_b8c7_1f1b_d998_9d07_c1f6;

        #200;
        key = 128'h8704_38e9_d311_48d1_175a_17f8_62ff_8f75;
        state = 128'hd0d4_f285_b109_32b0_a4db_b899_1a56_76ea;

        #200;
        key = 128'h95f0_0e00_4ae0_19df_ba15_d301_43dc_f5f2;
        state = 128'h0d4d_7a75_d5d0_90b3_e0ab_6a6a_77ce_9f11;

        #200;
        key = 128'h52d6_ed09_49a8_b972_91a6_1741_4c86_5e02;
        state = 128'h2f92_d713_1e1b_bcde_cc66_3383_8bf9_a2ee;

        #200;
        key = 128'h2109_a654_b46f_3f00_270b_0dd1_1f0f_8b33;
        state = 128'h9821_29b2_13df_9c53_bc84_5f88_fa4c_7daa;

        #200;
        key = 128'hb9e6_bb5e_cf88_4114_d0f2_1648_b503_fa5d;
        state = 128'hdd50_c9af_34f2_581e_cfb1_0a66_9801_c2a4;

        #200;
        key = 128'h7ed4_18f6_22b8_906e_8533_f6e4_b386_092d;
        state = 128'h5b70_a0d3_0570_05a9_7c21_3cec_d797_07d6;

        #200;
        key = 128'h426e_e550_8e1d_1be2_5284_2368_352a_532d;
        state = 128'h66d1_71c9_92f5_8b65_7951_58ad_ec30_b952;

        #200;
        key = 128'hab23_91bd_de18_22a4_ad54_f308_49e3_936c;
        state = 128'h144d_45dc_edf4_529c_2943_1e64_635a_7994;

        #200;
        key = 128'h4103_9883_950a_585e_54be_078c_4369_70e3;
        state = 128'h2679_7ff2_48a7_d641_7e87_df2c_1385_5153;

        #200;
        key = 128'hbba2_6704_ee7f_1bf8_07f1_0d02_8f6c_2762;
        state = 128'h663b_236e_b716_6cff_f793_f347_924b_c7f1;

        #200;
        key = 128'h3eda_dad8_500a_a746_c5ad_eff2_d623_35ff;
        state = 128'h4716_eac1_34a5_81ed_ca9f_0480_eec4_0951;

        #200;
        key = 128'h1753_41c3_be0c_ae77_4ff0_01b1_79a6_ee72;
        state = 128'h799e_04d9_2c9c_2dd5_125a_d0e7_c46b_914a;

        #200;
        key = 128'hd714_8c46_4b3d_382f_5110_6e2d_ccdf_027b;
        state = 128'h764d_af46_fefd_9cbb_a103_cd41_0228_5883;

        #200;
        key = 128'h37c9_32bf_ec96_809b_3269_cfd3_6026_3676;
        state = 128'h5489_29ab_6b30_4562_8d73_ee3b_0213_1c0e;

        #200;
        key = 128'ha9d9_58de_848b_d8ac_f888_43ec_814f_bc67;
        state = 128'h1f12_9e78_ce68_4fa3_907e_948d_bc62_2993;

        #200;
        key = 128'h8eb1_adc6_a548_be7a_04ee_eaba_4e46_68fd;
        state = 128'hdc25_eecc_df18_3742_d5c1_111b_1b4b_e2ee;

        #200;
        key = 128'h6bc7_fc8a_0cf6_4603_a5dd_cc3e_8e87_9037;
        state = 128'h880b_edd2_51ab_fce4_dd03_559f_c273_f9a7;

        #200;
        key = 128'h4d30_5185_2aac_9a49_6a4d_af50_94a8_6eab;
        state = 128'hc875_b1b9_2e07_5325_d8fa_f27e_51c1_f3ff;

        #200;
        key = 128'h4a30_7aa7_18bd_7109_cd1b_1969_6c32_7599;
        state = 128'h2d41_e301_39cf_15b4_7f65_7dc2_4e18_2198;

        #200;
        key = 128'h0703_b497_404a_b22c_6221_1938_a4df_7ca0;
        state = 128'h8855_6e6b_dce9_3c3e_7617_5463_33ae_ff69;

        #200;
        key = 128'h7a3d_58fd_1762_a192_e659_91fe_bbeb_4a93;
        state = 128'h52e0_a52d_86a2_d517_378c_b026_352d_9305;

        #200;
        key = 128'hc205_11a4_8aa2_ab03_ba7c_8e68_47dd_5a84;
        state = 128'h8565_7607_a67b_d8ad_98b9_fc29_4842_8202;

        #200;
        key = 128'hd88a_60f8_c18d_4ed2_588c_02cc_e61b_b1ad;
        state = 128'h67f0_bd74_0a2f_3fa6_7a00_7c1e_286d_e1eb;

        #200;
        key = 128'hbe7f_0176_28b5_3390_f309_1c03_6e68_116e;
        state = 128'h0c75_d150_50e3_b0a4_d059_5e8c_3b60_bc7f;

        #200;
        key = 128'h2cea_c1fc_2e16_5314_91da_6c2a_b274_23d9;
        state = 128'he844_cef4_3ea0_f207_4858_c332_c2a4_6c20;

        #200;
        key = 128'h80b6_f63d_b99b_83ef_eeb1_918b_8251_67e9;
        state = 128'hbb26_ac5f_dc23_9f04_a743_5fe5_9142_f40a;

        #200;
        key = 128'h0afd_ae91_3b5d_0008_5351_41aa_00d8_b524;
        state = 128'h217f_8b5e_2383_085d_ec35_2f55_aa98_e738;

        #200;
        key = 128'h9d7a_fe31_23ee_696f_75a4_ebe3_78e0_41f2;
        state = 128'hf8bd_289f_a407_0ee7_3b69_d89f_18d0_43de;

        #200;
        key = 128'hacd0_8466_0f83_6007_126a_642b_cfdc_5142;
        state = 128'hed25_d5b4_ae1f_12a4_bfbd_4438_54a9_1fea;

        #200;
        key = 128'h67ca_3cdf_5475_268c_8e16_39f1_d95c_7f27;
        state = 128'hcc2e_07fd_a81a_b3b3_6664_135a_78e0_c64b;

        #200;
        key = 128'ha28b_6afc_8957_b57c_58b9_926f_8e0e_3edc;
        state = 128'hc18e_87e8_d37e_f112_cdd5_59aa_4001_ebd7;

        #200;
        key = 128'h2d66_39e1_7357_8af3_6af5_41a0_dd00_710d;
        state = 128'hc29b_1f74_90f3_effc_db6a_cad9_1cbf_a33e;

        #200;
        key = 128'h85f0_1234_bad9_8095_c0a2_7284_1907_5b23;
        state = 128'h0388_10aa_14a4_44d9_3763_737d_378d_92b8;

        #200;
        key = 128'hc2f3_d26f_1c50_b725_4106_fbcb_e2c1_3ef2;
        state = 128'h00bd_e25d_eac9_66e6_a744_aca3_d021_4882;

        #200;
        key = 128'h50f4_edb0_61bc_aff7_84ad_6581_fbaf_b665;
        state = 128'h9cdc_fd96_d348_6158_85f9_af76_6255_62eb;

        #200;
        key = 128'h7679_5542_ca96_c407_b068_8034_acc3_c47c;
        state = 128'hbf00_9fb2_95ce_1d3b_fb92_90d4_d1f8_fd9c;

        #200;
        key = 128'h5185_f6dd_feb8_4dc6_ada8_ddb7_8c10_81a7;
        state = 128'h5761_9d73_1749_d733_b750_a3e0_7ccb_6a30;

        #200;
        key = 128'hcb15_c38c_de5a_ceb4_afda_8ace_6d4e_3181;
        state = 128'he012_e855_5cfb_9a8d_8b31_42dd_f701_03a8;

        #200;
        key = 128'hba74_cb42_1e2a_af90_a160_df23_c846_f3c8;
        state = 128'h1e84_60e9_9735_294f_3715_638d_2daf_0110;

        #200;
        key = 128'h5c9b_fabc_0a4a_b3a3_f545_1933_7ddf_bc2e;
        state = 128'h43cc_dbed_9a79_4d92_9513_9803_4b92_addc;

        #200;
        key = 128'h03b7_c104_f984_d2ef_eba8_f04a_001d_260b;
        state = 128'hd6a3_cb75_2fc1_4b82_f08e_c917_01fd_ec55;

        #200;
        key = 128'h1e28_064a_b8cf_d946_c50d_e72e_3533_ee09;
        state = 128'h6826_4d4b_8eec_9492_3488_bbf2_c470_9368;

        #200;
        key = 128'h0f08_23a8_5c2a_b9be_e33b_14f0_ab05_162c;
        state = 128'h8299_afed_6dbc_c9fe_238b_e150_ad15_1740;

        #200;
        key = 128'h646e_38d4_fab0_efa2_6f4d_aa30_e4d7_7027;
        state = 128'hfe21_ccd8_754b_d6bd_e142_ce91_58e0_9abd;

        #200;
        key = 128'h0d0c_d44c_43c2_be5e_224f_2e14_1dd6_8ac1;
        state = 128'h0a4c_81c7_33a6_c6fe_25d3_fb9f_8447_aa8c;

        #200;
        key = 128'hd51d_e3e3_bf2c_059f_c95d_16d0_f8b0_b8b5;
        state = 128'hcb21_e544_0346_ed31_f13e_7c8c_a152_2c81;

        #200;
        key = 128'hc470_2043_956d_73ec_00e0_bec5_20b8_81f5;
        state = 128'h3870_cd04_d245_0add_3c64_444d_e2ce_bdc5;

        #200;
        key = 128'h54e7_c9b4_8c16_0090_e3fa_7f25_c1a4_a44a;
        state = 128'h6c0d_e731_f5e2_98c1_8b56_adda_8575_bf0d;

        #200;
        key = 128'hadac_c080_fd33_d0f6_4655_30d7_de7c_48a3;
        state = 128'h1fc8_8ed7_c87b_3114_13c4_a7b8_fc79_e684;

        #200;
        key = 128'h1fc0_6480_43c7_9e9a_23d1_68d4_58f0_9f01;
        state = 128'h90fe_9931_193f_4dc2_11b9_2e1a_4dfd_6125;

        #200;
        key = 128'hee80_091d_d184_113a_dd70_7c51_0add_73ff;
        state = 128'hffe2_7475_f1a6_6770_f280_9b7a_75e1_cb50;

        #200;
        key = 128'hda4c_2e93_fc04_24f3_b93f_0647_4dcf_9b3d;
        state = 128'h860f_7337_55e2_74bb_18c7_a24a_3841_0eea;

        #200;
        key = 128'hb08c_a7a8_ff46_9a47_9c2f_1052_ac9a_f2f4;
        state = 128'h827f_07b7_5194_a0e7_8ef1_fecd_e209_29af;

        #200;
        key = 128'h49ed_c6e4_1858_f163_2a20_64f3_a004_85f7;
        state = 128'h14a7_81e4_1244_e941_01be_661f_c953_5232;

        #200;
        key = 128'h9354_d1cf_be64_8874_47dd_384a_13e0_2b0c;
        state = 128'hd012_4064_404b_d6df_dbc5_76d6_ad5a_507c;

        #200;
        key = 128'h3165_628f_9d53_6067_033b_ff63_6eb7_1d2f;
        state = 128'h9a94_ca13_e1f3_1072_1e34_a7e2_35b9_d3f7;

        #200;
        key = 128'h646b_eb1c_e30d_744b_89e3_268f_7106_ad83;
        state = 128'hac36_aa9b_74f5_f69d_753f_4d3e_7ef0_f70b;

        #200;
        key = 128'h5ee0_eccc_c1ae_178b_690c_2050_0841_87f2;
        state = 128'h3799_c02b_8063_560c_0fe2_017c_770c_471f;

        #200;
        key = 128'hd12e_8b8f_7b2b_4533_a5a1_f050_bc5e_2d28;
        state = 128'hd81d_05f1_4b05_1005_fae7_a51b_96ff_5629;

        #200;
        key = 128'h63aa_d7c5_af3a_9a2a_af0a_3715_ac6a_53be;
        state = 128'hebfa_4c9d_79ca_5379_ebfe_1709_01a6_5977;

        #200;
        key = 128'h8609_bd4a_d2da_40cb_c4a8_af7a_754f_f005;
        state = 128'hbaf3_b6ba_a4c2_f760_cb54_948b_8635_df57;

        #200;
        key = 128'he5de_e1db_c7db_45b0_aa77_b2d9_d2ef_b2d0;
        state = 128'h0b5a_0a4f_f2ab_9bba_de24_cd32_1377_8a8b;

        #200;
        key = 128'h1c21_ab7e_7a10_5fe5_86e4_a974_3efd_6b64;
        state = 128'hfd48_a2df_ccd9_827d_385b_a5c2_e5b4_1bc3;

        #200;
        key = 128'ha7da_3cb7_667c_6f9b_3ca2_fc58_3563_1fd4;
        state = 128'h7bb1_a665_485e_59f2_646f_dee9_5f6f_f657;

        #200;
        key = 128'hba91_17cd_6c3d_4397_0be6_0594_30a6_6d2c;
        state = 128'h3dcf_f824_7b3e_b34b_369d_be49_d08c_789b;

        #200;
        key = 128'h3b1c_59ca_71df_ae29_71bc_79a7_313f_793c;
        state = 128'h5ecc_333b_b000_4c15_a919_1f17_1585_34cc;

        #200;
        key = 128'hd4f7_94e4_bc92_f2ce_c8bb_7e4d_3a02_094a;
        state = 128'h0392_9276_f52d_4bc0_fbe3_d8b9_5da9_6174;

        #200;
        key = 128'h544a_32b0_4281_a587_80d3_deb1_8313_6a18;
        state = 128'h7f5e_80ce_206e_bfe8_076c_a0f8_83d0_9244;

        #200;
        key = 128'h6fb5_7ec7_67d2_a5ca_064f_e698_1d07_b7b6;
        state = 128'hb01c_8e94_b5d3_6808_a93b_74fd_5bc2_1b65;

        #200;
        key = 128'h02ac_51b4_a6cd_05ce_85b2_3d1d_a2cb_af9c;
        state = 128'h3212_c2a4_4492_c3d2_9955_dd24_620a_8f72;

        #200;
        key = 128'haf14_494e_23ae_d865_f2cf_2b46_a067_cc1a;
        state = 128'h66a6_9a8a_ee4b_5776_9544_9c1b_3bb2_db96;

        #200;
        key = 128'hd368_ab21_585c_313d_2175_78dd_5fc8_4429;
        state = 128'hc443_b679_0bcb_d5b3_4243_7a0e_93c3_6781;

        #200;
        key = 128'h3215_a452_886c_d6da_4be4_250a_6aa8_e24d;
        state = 128'h55a6_ec40_e489_26a7_4f09_3863_284f_4179;

        #200;
        key = 128'hfd3b_49a5_f14b_847d_0728_c131_47b4_7480;
        state = 128'h671c_080b_db9b_c46d_077e_6354_1cd5_9794;

        #200;
        key = 128'he462_6b4f_408a_9564_732a_5749_88f6_ff7e;
        state = 128'he8cf_d7e2_e174_0adb_ca71_8045_571f_6f04;

        #200;
        key = 128'he70f_f4a2_e3ca_1c1f_f00f_81de_31af_9447;
        state = 128'heee9_d556_5577_7776_eef2_0cf6_1a2c_4a55;

        #200;
        key = 128'h4aff_a705_910b_8933_6688_9889_c2ec_bf1d;
        state = 128'h7698_cdb0_41ea_313e_74dc_06e1_b0c6_da85;

        #200;
        key = 128'hc485_abf0_1563_5340_1176_2c30_790c_de7f;
        state = 128'h3729_49ea_a486_a5a6_2dc1_082e_c2c7_07a3;

        #200;
        key = 128'h4caa_5434_d516_50f7_f618_c1fd_e4c5_6615;
        state = 128'h3f64_864e_6723_735e_8e62_0eed_b32d_e434;

        #200;
        key = 128'h437b_3250_0874_ec65_dde8_6f15_2d02_1246;
        state = 128'hfade_5581_8964_d22d_2e22_a917_dc0e_37b1;

        #200;
        key = 128'h4ddc_f4e8_09fc_6d16_ee88_23b8_dd1b_ffd8;
        state = 128'hfe0d_130f_e007_287c_ce7b_ceb8_f8a9_bd56;

        #200;
        key = 128'h48fc_c081_d3dd_773c_3c38_40c0_526f_e69e;
        state = 128'hfb72_144a_b078_ca8f_8d75_e556_7209_5550;

        #200;
        key = 128'heb2f_a8f9_6b77_c68a_4231_febd_77d2_4538;
        state = 128'hd20b_5364_0473_d980_e2c1_039b_d965_4082;

        #200;
        key = 128'h28e9_055c_6168_5ec5_ab02_f362_e11e_b235;
        state = 128'h77a6_9b3a_e05d_e1ac_a212_dac6_99ee_14d5;

        #200;
        key = 128'h710f_ec7c_1a09_3445_519f_58e2_8d39_9aaf;
        state = 128'h38a7_c384_fcbf_42d7_205b_5d9e_e8b6_8d7c;

        #200;
        key = 128'h23c5_e3f5_bfea_d7d9_1959_ac0f_0407_10df;
        state = 128'h2a9d_228d_73d5_2023_d5fc_b228_4a67_9d54;

        #200;
        key = 128'hc58e_85f2_04bc_8078_783a_260b_0463_3ede;
        state = 128'hed07_d1e0_0929_fe8e_d7b6_1df0_117d_99b0;

        #200;
        key = 128'hc692_1aa8_dbfa_f11a_3a3a_68bf_180a_beb6;
        state = 128'h1861_ac1b_9b36_2ba4_0f25_5051_5255_88a1;

        #200;
        key = 128'h60f2_02f1_2adc_d5eb_5649_0fdf_488f_38d7;
        state = 128'hb294_9655_b4b2_a6cd_2b74_1fc5_90ee_b2ef;

        #200;
        key = 128'h3e4c_5b42_1f4d_0144_3b1e_402c_0250_2190;
        state = 128'h64ff_32bb_105c_253f_107f_6048_bf8e_d6fd;

        #200;
        key = 128'h2a3f_febb_9a38_f86e_fae5_8e55_5e7d_c809;
        state = 128'h43bb_f690_68f3_51b8_c483_bcd8_b97f_2ee8;

        #200;
        key = 128'h2841_e362_d1ef_5981_bdc4_f5e6_53bc_abd4;
        state = 128'hc8a7_a13b_9120_a416_d49b_f433_3b1e_9868;

        #200;
        key = 128'hd467_8a4d_def3_8e17_894a_611c_4586_0915;
        state = 128'hcf15_5253_4bb6_b60e_ae2c_f0b5_67cb_ac39;

        #200;
        key = 128'he88f_379a_1f69_58be_632e_cabc_8a7d_882b;
        state = 128'h0db8_0d1f_cafd_ac1f_d097_30d9_f032_39a3;

        #200;
        key = 128'hb5a9_b433_1a87_a210_179a_6b44_4cf2_3c87;
        state = 128'h72ea_84ee_6cb1_0cfe_255f_a300_1fda_b56b;

        #200;
        key = 128'h112b_a4eb_a9e0_f45a_8f9f_689a_b7b5_730a;
        state = 128'h8844_a784_06ca_a92f_8aee_8393_db29_b3cb;

        #200;
        key = 128'h57bb_7de2_54be_4b1a_c417_5c7f_4b6a_0284;
        state = 128'he068_cff0_96a2_817e_bed4_af98_1800_e0c0;

        #200;
        key = 128'h82a1_82bb_a81c_7211_c9ca_bcc0_9567_5fc1;
        state = 128'h590e_a1bb_c0a2_6ad1_1f01_f2de_a6cb_68b5;

        #200;
        key = 128'h78eb_e99c_7a51_71ef_4090_17ef_8e59_c451;
        state = 128'h0d15_879f_e0a4_867e_53ee_af09_3926_6fff;

        #200;
        key = 128'h645d_0acb_3f71_f08a_9bea_e69f_7992_62d7;
        state = 128'h8fc8_b0ce_ebe4_5ea6_88ea_3739_7503_276b;

        #200;
        key = 128'h6bd0_93cb_2bc6_8edc_c30c_4f9d_f4f3_2a30;
        state = 128'h8673_05d3_8dfd_bdd5_55e3_fb4d_5a05_e30b;

        #200;
        key = 128'hf53f_1050_30dc_7c90_90d0_db8b_0490_08a1;
        state = 128'hf070_2ea1_438b_b9ce_bebb_6a86_fb85_7298;

        #200;
        key = 128'h1a61_c78c_4252_2cd6_9425_dbdc_f87b_b3d0;
        state = 128'h4c8d_da34_85af_1699_bfd8_edb1_f325_15d4;

        #200;
        key = 128'h61d8_e40f_2c87_06de_2ac4_b2b3_d18b_dbed;
        state = 128'h48c8_26e1_ab6c_30c6_7e3a_30aa_95d4_961d;

        #200;
        key = 128'h3ff7_72d7_ba60_195f_198b_4aaf_40d6_a8f4;
        state = 128'hfc1a_4753_a6f6_b71d_fca3_3f67_09f1_a8f5;

        #200;
        key = 128'hc510_4bbf_f222_4aad_4bb2_66c4_4b10_02e9;
        state = 128'h0e16_0d35_9b9a_a962_7764_743b_fa75_f831;

        #200;
        key = 128'h2704_bb90_5246_01c4_f2fe_710b_8d65_5d63;
        state = 128'hd161_5333_652f_cf79_35b0_5e23_19cb_8a0a;

        #200;
        key = 128'h2464_0b78_8635_7ecc_6cf7_3229_54cf_3fc5;
        state = 128'h2ca1_ca2c_ba41_a963_b9b7_0e0e_b88a_ff1b;

        #200;
        key = 128'haa66_01b8_6c04_b88e_c47e_36e4_15c9_86e1;
        state = 128'h582b_1793_3aab_51da_ac4b_3b63_be09_ef0d;

        #200;
        key = 128'hbbd0_591f_e1e8_de3f_2c69_8d42_e8ce_e474;
        state = 128'h3080_db24_bb2b_d470_0394_4ab8_9e2b_ef7c;

        #200;
        key = 128'hb3e2_0ad6_ed28_16fe_c0fb_9be1_5afb_6f5d;
        state = 128'he176_0a14_65df_2616_bdc2_1830_63e3_5f61;

        #200;
        key = 128'he0c9_5df6_a636_962b_c4c5_e125_5e89_f2e8;
        state = 128'h99d1_d6f3_6c8c_dff8_4056_399f_c21c_454f;

        #200;
        key = 128'hee49_1183_602c_9083_2d17_3c66_9475_fb4a;
        state = 128'h741f_7ca1_c32f_20dd_8617_bd65_23af_4928;

        #200;
        key = 128'h0579_19a1_4d16_179b_f0a1_0f39_940f_0f3f;
        state = 128'hbd63_42d5_1821_d219_1a1e_daeb_a14e_088e;

        #200;
        key = 128'hf69f_0f2c_4945_336d_dea8_f282_b658_f43d;
        state = 128'hdd4c_3140_2090_8ee7_7e3e_76f4_4bbb_b99e;

        #200;
        key = 128'h86a3_5be9_57b6_92f1_82f8_0cdc_9b60_8e55;
        state = 128'h5c65_683f_a0fa_eaca_b081_1b7d_5799_e718;

        #200;
        key = 128'h2dce_9c7f_2580_2915_7019_f2bc_6872_b743;
        state = 128'ha9d1_a072_604a_1505_151f_facf_bc5a_4c9e;

        #200;
        key = 128'h8e8c_3ef3_ad2d_bb3f_4edb_7a17_098b_7581;
        state = 128'hb408_d344_d5b0_8bc7_caea_a5e8_524f_33d9;

        #200;
        key = 128'hfc22_225a_36c4_47c0_e27a_5102_b282_0352;
        state = 128'h4ddb_59d6_04d4_a8af_e24e_5c12_bd65_bac9;

        #200;
        key = 128'ha0c2_6b12_f300_9253_21f3_be96_8b95_6bd8;
        state = 128'hc016_c431_f3c5_89a6_04d8_e26d_53e7_0fc7;

        #200;
        key = 128'h7b86_22c7_d120_78d9_4b46_45a9_5c58_63ef;
        state = 128'hed2f_bb20_ff84_76c9_099f_0086_02b0_a46b;

        #200;
        key = 128'h05fe_b95f_6815_4518_da5c_aacc_246f_7757;
        state = 128'h681d_351c_7529_bb7b_312c_1710_0352_0d26;

        #200;
        key = 128'hbef4_a4cc_797b_26e1_6933_ddbb_87c6_8216;
        state = 128'h31ad_a932_eda3_03c9_e4ad_0a31_0607_fe01;

        #200;
        key = 128'hf311_3a01_9cee_a509_8a59_1adf_8b0b_a052;
        state = 128'h90a5_5315_d135_8781_68b0_2a10_2011_e485;

        #200;
        key = 128'ha4d7_a342_f258_abce_b794_0255_2bbc_c906;
        state = 128'h6922_e468_16a0_7cf3_c4f3_4af7_0d9e_843c;

        #200;
        key = 128'h3a75_2bb1_c1a1_386d_7bd1_2967_96c8_15af;
        state = 128'h90ea_2580_1709_77e3_91af_a9f3_1bac_6735;

        #200;
        key = 128'h3379_867e_4c8b_bf9e_8567_4049_6308_9be8;
        state = 128'hbb81_4f4f_2208_96ae_5bff_ec90_d966_2db9;

        #200;
        key = 128'h7a4b_6f7d_bb0a_9230_21a4_664f_3bcb_5f0d;
        state = 128'he55c_3085_c098_ff60_ae81_c234_55b5_e55e;

        #200;
        key = 128'hff12_3341_848d_395a_b699_9b7f_d425_25a3;
        state = 128'h51b3_382b_299c_9fb2_28d7_79e6_c05c_583e;

        #200;
        key = 128'hd5df_8c95_9f99_96e6_f31b_ac71_50bc_8f3d;
        state = 128'h2775_84cb_8266_b45b_2d07_153a_36e9_59d6;

        #200;
        key = 128'h9689_c98c_2d97_f0f1_0236_47d7_57eb_90d1;
        state = 128'hb08f_0010_d710_28a2_2ba2_fb1d_559f_2371;

        #200;
        key = 128'h1a9a_517a_b19b_3b51_6d57_d556_613f_2375;
        state = 128'h5ba4_2da2_f88d_0b84_14c8_5041_3aad_2e02;

        #200;
        key = 128'hcfdd_5e97_59fa_0a46_d986_a88a_1a9e_d428;
        state = 128'ha83e_ec64_4418_3aa1_1617_90ef_de5d_fc31;

        #200;
        key = 128'h2a5e_ddf0_fbba_7980_9078_76e4_bc35_b689;
        state = 128'h5f70_9769_3319_a419_d516_b3a5_d493_8342;

        #200;
        key = 128'h205c_ebf7_cc5a_25f5_951f_41bc_522b_1f92;
        state = 128'h6061_6369_2319_f258_7dc1_9e78_19b1_a012;

        #200;
        key = 128'h9064_785e_85bc_03b2_20d4_0556_e211_bf14;
        state = 128'h9be7_3e72_74a0_582a_3faa_5054_8bab_786d;

        #200;
        key = 128'hf7ae_8d6f_f677_f7c9_6622_b2e2_58d7_2866;
        state = 128'h0698_b68f_2316_71f9_aeb0_277a_fdb9_e430;

        #200;
        key = 128'h586c_4b64_79d5_9e6d_f78e_9704_2ac7_ee33;
        state = 128'hf6ec_38e6_73db_3e46_af8a_3dad_b25c_bbb4;

        #200;
        key = 128'h6c05_bc0c_0f98_065d_ec7a_4501_466a_dc50;
        state = 128'hb3f4_9a96_889a_e1cd_5d87_f4f9_dd09_9039;

        #200;
        key = 128'hdc5a_448c_2f94_b3ff_80a7_7395_8ba0_bbe2;
        state = 128'h4597_1edb_4143_adff_8436_e4b1_aedd_9348;

        #200;
        key = 128'h0c3b_9ae2_4be0_d05e_8c7e_d7f3_45ad_8079;
        state = 128'hd599_a310_86fd_507f_5a74_cc87_f848_e7c6;

        #200;
        key = 128'h3879_1d58_5bae_2577_4725_a06c_72bb_fe01;
        state = 128'h405a_31b4_d82a_fbc4_599c_d32d_ab0a_ec8d;

        #200;
        key = 128'h5729_1e8e_ea73_8887_7814_332a_4576_f0c7;
        state = 128'h1ca6_3af1_9a0f_c966_023e_9b87_6714_230d;

        #200;
        key = 128'hd424_1c6d_f3ea_0172_843d_65a2_e633_b303;
        state = 128'hfc5a_fb79_eab0_00d6_1759_5373_8317_54ec;

        #200;
        key = 128'hb0a6_0860_a044_d047_5e5b_1258_8bb5_c2bc;
        state = 128'h5765_d53f_68c9_5c1a_f964_4474_c7f6_ce79;

        #200;
        key = 128'hfe54_f510_c7dd_9fa2_d069_7e17_bf38_c487;
        state = 128'h1e70_e862_968c_9044_1e1e_ef62_a0a8_463a;

        #200;
        key = 128'h3b1c_7de1_7f60_f4f3_ca85_70c3_05e4_a6f8;
        state = 128'h2e1c_aad8_8b63_7123_a3ba_ca87_ed0f_8dd1;

        #200;
        key = 128'h0e33_4cae_d9b5_6822_c9ef_f594_92b9_8da0;
        state = 128'h35f2_dcd5_1967_71ad_6b57_8c0f_19f4_9811;

        #200;
        key = 128'h4f87_f0e8_a1ad_de01_ebf9_a072_7706_83e0;
        state = 128'h4352_6825_1c68_727a_3171_82d7_f04c_40d9;

        #200;
        key = 128'h4d13_a439_3687_9cfa_b8b3_491e_b365_f249;
        state = 128'hed05_5328_f473_1e7b_48e0_23c3_afe7_2cee;

        #200;
        key = 128'h283b_5653_c2fb_289c_3263_48ec_2349_fb04;
        state = 128'h29f0_0082_b8ea_cbb1_f0c7_0d70_31ec_a673;

        #200;
        key = 128'h610a_e261_88dd_f3d5_ab06_d6fc_ef23_9189;
        state = 128'hbe0f_ac89_99eb_e146_2356_566c_a06b_ad7d;

        #200;
        key = 128'h3f2b_1425_6159_0f45_3a4c_db1b_c106_acc7;
        state = 128'h5d09_c908_b48a_25a5_7a8d_9c02_218e_085f;

        #200;
        key = 128'h2e79_8cbf_c721_a7e1_81b9_7aaf_2956_a958;
        state = 128'hed89_d99c_b8f1_7764_d299_2676_bc5d_67b1;

        #200;
        key = 128'h9b0b_4249_80a2_cb8e_0a5e_1377_6fe4_1724;
        state = 128'h50dd_9479_ab58_3be6_aa1f_0bdd_b6ec_8bb6;

        #200;
        key = 128'h9a0c_1cef_ba68_f678_e164_96af_53da_595b;
        state = 128'h975e_586f_200f_c75d_8fc5_e34d_5c75_9b78;

        #200;
        key = 128'haa02_7a88_a759_f058_4eca_da3b_1e23_fcbd;
        state = 128'heea1_704d_f318_b4f6_d20a_9171_5f6f_c542;

        #200;
        key = 128'h1cb0_b540_f393_20e7_2e7e_5033_ad92_ef43;
        state = 128'h3995_5288_35d6_672d_cf77_d77f_1bf5_d722;

        #200;
        key = 128'h9a58_1470_3899_7cab_a6b5_4856_e955_1d54;
        state = 128'hde07_0097_b4f6_5e35_396d_0a8c_377d_73d9;

        #200;
        key = 128'hdafa_c7a7_7292_d640_ddf7_d32f_a23e_a934;
        state = 128'hc5e1_90cc_9817_bd30_4a67_2e17_dbda_60ca;

        #200;
        key = 128'hbbf2_c314_8638_d720_e8f3_e518_b309_d0ed;
        state = 128'h8f2a_c63a_ea06_ab98_5fe4_676a_64c3_85f8;

        #200;
        key = 128'h6584_fe9c_fe75_4b6c_b98d_fefb_f878_539b;
        state = 128'h9592_9a3e_4f4d_e3ec_be7d_160e_704e_e60b;

        #200;
        key = 128'h2bde_7987_544d_b0fc_4b7e_e8ea_de7e_26f1;
        state = 128'h6ce8_2ea4_e29d_f206_b926_6d5f_fbbd_1739;

        #200;
        key = 128'h8659_d4b4_570f_253d_3344_84f4_cd35_e108;
        state = 128'h5957_742e_87cc_6554_3a88_d560_c375_3432;

        #200;
        key = 128'h4c96_9b4a_d84e_c136_be81_a469_c504_e9aa;
        state = 128'h1fcf_e8ad_485d_d142_722a_9eeb_cf25_d5d7;

        #200;
        key = 128'hc0e0_f976_f993_1ca7_8232_0fa2_f602_a0a3;
        state = 128'h6f63_8eca_e8e2_4b8d_9c57_8de2_a772_bb8f;

        #200;
        key = 128'h67df_491a_d557_08f8_dbc9_2290_d27a_4fde;
        state = 128'h50ee_8faf_cff0_f000_0926_e41a_fb1f_27f9;

        #200;
        key = 128'hc612_f59d_de67_60a1_30b8_db7c_7ed4_e56a;
        state = 128'h21df_db30_c020_09ba_757c_1f97_f15e_0a80;

        #200;
        key = 128'h85f4_fe78_d0c9_0a37_fbba_da21_9a47_4010;
        state = 128'h2b4f_dd1a_55aa_a7ab_bf56_a6dc_2b15_a1b9;

        #200;
        key = 128'h4a2c_4982_b80b_8057_32d4_2606_8ad6_ec6c;
        state = 128'hddd0_a123_94e2_f0ee_e3d0_796b_4ab4_bac2;

        #200;
        key = 128'h61f4_d90d_fe2f_718b_9c89_695c_4ee0_12d1;
        state = 128'h4ea8_1abf_1f2e_6b10_2ed4_8bf3_92ce_eaf7;

        #200;
        key = 128'h5f40_dc14_1d27_4851_b478_f451_caeb_e051;
        state = 128'h682a_0797_4f05_7d2d_6dd6_753c_f9fa_cd69;

        #200;
        key = 128'h5e0f_86fa_39af_71e1_7865_a4e1_fdf0_967f;
        state = 128'h2b69_988d_5390_6e45_aa7c_598f_1a1d_e23c;

        #200;
        key = 128'h23a5_7fb3_d349_3d66_c9e2_cbbb_1378_7fd9;
        state = 128'h0c4b_cc9d_c325_0b03_01a8_76f8_f29f_19fb;

        #200;
        key = 128'h57f7_5c03_dfff_f8c3_5f4a_7d52_7cad_d208;
        state = 128'hd4dc_4367_df54_53f3_32ac_f5db_cf06_d508;

        #200;
        key = 128'h3c39_228c_2856_2b9c_7724_927a_e01f_7a25;
        state = 128'h4159_a354_5a72_16ae_6c27_a1cd_89ec_0b7d;

        #200;
        key = 128'h98ef_b7e7_b620_87c2_4127_2d84_1a87_a58f;
        state = 128'h5287_945f_b20e_2b3a_4f30_2965_97cb_43f5;

        #200;
        key = 128'hb13f_32ef_6f47_a2cc_9c4c_928d_be08_2dab;
        state = 128'h3b71_6555_e515_7606_c5ba_2fed_4e42_c566;

        #200;
        key = 128'hcb54_2160_46eb_1084_c52a_3afc_5c60_8ddd;
        state = 128'he3df_0f2e_5f2e_8e74_b7ef_0980_d2f9_5524;

        #200;
        key = 128'hdb5e_8fd9_9409_309a_afc8_4d67_de6f_5abe;
        state = 128'h2d05_12f3_2083_4173_b32a_8278_b302_de13;

        #200;
        key = 128'hc086_08ca_c061_d562_c9c4_4283_5d77_07db;
        state = 128'he39e_9b20_ef61_dfe1_b3f8_8046_a05c_a9c9;

        #200;
        key = 128'h0ede_4d69_402c_10d9_7811_64d4_7e7b_dbb0;
        state = 128'h9fba_ee2d_ea71_dba5_56e9_d011_0433_abf0;

        #200;
        key = 128'h7900_2acb_b472_b97e_c7eb_356b_cfeb_0fe3;
        state = 128'h9a72_1474_0a65_485e_1600_6659_09e6_1c4b;

        #200;
        key = 128'h6501_00ed_d936_4ec4_66e5_c38b_ae10_30cd;
        state = 128'hf70c_fee6_9e3a_5a90_764f_4e5a_e4cd_cd60;

        #200;
        key = 128'h2ace_c706_f17f_e039_c5c2_3e83_2164_4206;
        state = 128'h40a6_893f_f81a_e92b_2d1c_89b6_af2a_ec05;

        #200;
        key = 128'hb9a3_052a_058e_b251_24a8_1905_da55_af22;
        state = 128'h3ce3_7bdd_b26e_2ec1_d38f_93b9_26d9_90b4;

        #200;
        key = 128'h1834_5942_9b38_8019_43da_22a3_713e_0a9f;
        state = 128'hc93d_f7f4_f323_0a92_b162_6fe3_2750_0ee2;

        #200;
        key = 128'h2f75_61b2_41e5_9279_5758_d73f_27cd_b2d0;
        state = 128'h5c17_5c99_a441_5e88_110f_cd39_5632_cc4f;

        #200;
        key = 128'h5cd9_f5f4_3e2e_46f1_16d4_d58c_bd09_8328;
        state = 128'h02f9_ecae_4fb2_c21d_99ee_7fa6_ab77_fcf2;

        #200;
        key = 128'ha094_5b1d_fdaf_7d59_5421_43b9_e05c_1cb7;
        state = 128'hcfe3_9f82_4b1b_24ab_bde8_9216_a03d_01a1;

        #200;
        key = 128'h5c4c_d771_7b8b_7a0f_3d35_4285_27c1_13b2;
        state = 128'hf1d1_7bae_5500_32be_1777_d093_edd0_a2aa;

        #200;
        key = 128'hb2c2_bf10_6b60_831e_3172_0cbb_7062_3b3f;
        state = 128'hfe6b_f7dc_ce8e_8beb_a3bd_a0a2_1ef7_f05c;

        #200;
        key = 128'hccd2_1635_2931_76df_d4c2_0cc2_e23a_094b;
        state = 128'h35d3_3f35_34f6_f216_39ef_9d79_08a9_9d9f;

        #200;
        key = 128'h305a_c08e_b0b2_9ec9_a8cf_9b75_92a6_ffce;
        state = 128'hc87f_47d5_2f73_ec58_23f4_de28_8d18_d254;

        #200;
        key = 128'hd612_72d8_deba_bfb5_440b_0b29_3a7d_e7f8;
        state = 128'h0428_55a3_2968_19c8_5544_f1c1_2a7e_2933;

        #200;
        key = 128'h8aa9_876c_7632_b6d4_368d_2ccb_9a74_5dc6;
        state = 128'h84bb_331c_1901_074f_40df_f18c_63fa_b2bf;

        #200;
        key = 128'h0558_6f42_f69a_9baf_4a3d_1157_dbed_c3df;
        state = 128'he325_7b20_f83c_650d_18fe_0695_1ca3_cf6c;

        #200;
        key = 128'h87bd_8a7d_433c_5328_266c_4817_7263_b9fb;
        state = 128'h0e32_fa2b_299f_0c41_a99f_8f3d_11f3_3ed0;

        #200;
        key = 128'hbf59_032e_b870_e66a_7f8c_8349_2418_3b0f;
        state = 128'h31ee_025d_5c7b_c3cf_0bd3_499c_42c3_8dca;

        #200;
        key = 128'h4ddf_5a3c_37d3_8534_5531_0144_2dd5_25ee;
        state = 128'hf5d8_9e29_a27e_198e_0a75_1495_1c10_f5a2;

        #200;
        key = 128'hf19c_e349_80a9_dae6_a039_2c70_6d60_752a;
        state = 128'h064b_74f3_8716_2a95_ddae_aa32_c5b2_48da;

        #200;
        key = 128'h9dd8_7a87_26e6_1503_d9eb_6513_45fd_2d3f;
        state = 128'hbdd4_efe3_3f8c_270d_73f2_80c8_7e98_1836;

        #200;
        key = 128'hed54_260a_903e_5745_e5e6_05dc_9d29_5037;
        state = 128'h2552_acd2_d5fe_b348_ad36_6086_b7e2_91f2;

        #200;
        key = 128'h7ab3_8a81_b26a_980d_01f0_1020_9cf8_0728;
        state = 128'hdc8f_c241_a4ac_c36c_b370_340a_df9d_7fa3;

        #200;
        key = 128'hbf23_de77_d938_860a_652f_d675_6372_3901;
        state = 128'hb6d2_46f6_99c0_a0f7_4fd5_8a51_140b_a025;

        #200;
        key = 128'h97cf_276e_0fbc_e4c1_c57f_aaec_41bd_3fab;
        state = 128'h7e11_6534_657c_9c89_93d5_9ff1_a9bf_8775;

        #200;
        key = 128'hf249_8a55_7601_58c2_fcd7_2502_fff8_a56c;
        state = 128'h6667_f13e_f33b_5a7e_c988_21e8_96aa_80cc;

        #200;
        key = 128'hc494_155f_25e7_8b2d_1316_1c94_7880_1343;
        state = 128'h4d0e_cbe4_08fb_35b7_cf14_6a33_b7a3_a41e;

        #200;
        key = 128'hc819_8828_4150_1489_933c_cf39_fc95_4af9;
        state = 128'hcdeb_2d91_b913_9030_afec_8403_3ef8_a824;

        #200;
        key = 128'h9c83_5a69_e7fd_3396_f974_3a97_131c_62db;
        state = 128'h2e6f_4610_436d_f7ea_90be_a18f_70fe_fb68;

        #200;
        key = 128'haf8a_5286_b9b3_c6a6_0e55_8ebe_7f93_47e3;
        state = 128'h9417_0023_3259_7950_aca2_fc02_f8d0_0df7;

        #200;
        key = 128'h970e_d557_e90b_fd03_0ce0_8c34_cb67_c992;
        state = 128'hd3ea_e237_6a18_601d_d149_8972_3704_198b;

        #200;
        key = 128'h289b_a7ef_a994_dcf7_c49c_0b3d_0364_bf1b;
        state = 128'hee65_3d40_e268_091d_0b75_907c_5691_2b66;

        #200;
        key = 128'h42dd_44c0_bb60_8eb6_4b32_6e4d_5e20_2605;
        state = 128'h15d6_3469_ee73_8035_e662_98d8_bd5d_27da;

        #200;
        key = 128'h57f1_5dda_1dc4_8a22_64c6_a6b3_e0ee_0302;
        state = 128'h5447_3840_0078_3d9f_76c0_1765_0c2c_7649;

        #200;
        key = 128'hcd41_80fc_fc74_7fa4_5559_6304_c6a4_137b;
        state = 128'hec8a_aefc_ea8b_c804_3b60_e062_b418_3d12;

        #200;
        key = 128'h33a2_76ae_4ba0_7720_74ff_a9f3_aa1c_be67;
        state = 128'h0f22_8d9c_ec84_d65e_ce6f_3d16_da36_21d2;

        #200;
        key = 128'h2c65_bf6e_c2ee_65fa_5c04_6725_3199_be5f;
        state = 128'h22a2_5247_5ba7_c8a1_632c_39fd_6949_b62c;

        #200;
        key = 128'he3b6_d7a3_7dd2_299e_c601_177f_4b53_4c60;
        state = 128'hf44b_d6e0_d016_6f56_b5ea_324f_0c71_71a9;

        #200;
        key = 128'hf594_bf90_4b31_40b7_f290_0cf5_388c_88a4;
        state = 128'h1215_1967_75d0_c0c1_e339_e5e5_6a31_887e;

        #200;
        key = 128'h73e3_9998_1310_1c10_9b99_3699_4389_7c84;
        state = 128'h12b1_98fe_f0af_5467_712d_a1eb_ef37_8d24;

        #200;
        key = 128'h7a86_6ba4_fd72_7f6e_6a07_7a7a_9c70_7423;
        state = 128'hb706_3aec_848a_f3a1_67da_530a_b870_20a5;

        #200;
        key = 128'h801a_9ad8_6c7a_db93_91de_ece9_bf82_31cd;
        state = 128'he61a_9026_abd5_19f7_b865_4b2c_d817_8f7a;

        #200;
        key = 128'hc86b_9e0a_0d96_7471_0d12_d416_e108_8a3d;
        state = 128'h6a5e_df0c_844d_7d60_f003_0ad6_bbcf_2df7;

        #200;
        key = 128'h4a6d_e9d7_b792_23a6_0556_be0f_b974_8423;
        state = 128'he750_9e2a_24bd_6388_a81e_4533_e523_840f;

        #200;
        key = 128'hd379_ff92_da20_30af_a29c_6ab3_dbcf_630b;
        state = 128'h483b_be3f_0855_01c8_374f_3a13_d592_1aa0;

        #200;
        key = 128'hdba0_2ce1_957f_ec4d_dff7_770c_7ade_cf44;
        state = 128'h28f3_4472_7cad_d691_5479_99ed_290c_fb87;

        #200;
        key = 128'h0d6b_c2a4_232e_8a1d_6577_fedf_9164_2b37;
        state = 128'h8227_b55e_6ab4_c987_cb37_3f83_9f86_2b0f;

        #200;
        key = 128'h2c86_7251_2021_04f8_7ef3_ef40_fc6d_981c;
        state = 128'h53cc_348d_15a3_24b7_6989_0007_4d5c_b913;

        #200;
        key = 128'h965c_afe0_fb6d_070f_6726_ba2e_e598_0c20;
        state = 128'h7564_4c44_1601_889f_c129_fd80_d945_c848;

        #200;
        key = 128'h9388_115b_d799_b821_c3da_ef47_acac_f57e;
        state = 128'hf52f_60c1_eb89_ab42_0be1_5f43_cb84_d5d4;

        #200;
        key = 128'h2ff5_29da_0863_bc12_5eef_e336_d1e3_c8f4;
        state = 128'hd2ee_175b_e6e3_46c0_058c_7469_80d1_0ec8;

        #200;
        key = 128'h9321_e23f_8614_069e_7f19_9552_3f2e_58c4;
        state = 128'h518b_16a7_1feb_6c2f_894b_bc03_2ff3_1d96;

        #200;
        key = 128'hfd60_6647_872c_4669_37fc_9bbb_6865_2354;
        state = 128'h807e_8601_01e4_d3e5_228c_4005_a080_379f;

        #200;
        key = 128'h13f6_eb88_cb87_b7f9_1061_273f_891b_6c99;
        state = 128'h7542_07da_43a4_9dd5_33a9_f711_60e4_769f;

        #200;
        key = 128'hc065_75d4_0cfa_14a1_12ca_4c87_d6b9_2e90;
        state = 128'h6358_ea79_f2e8_91cb_d0d4_2bde_cb36_f785;

        #200;
        key = 128'h4594_f407_6eee_2299_357d_8f05_2f90_00ac;
        state = 128'h96c6_696f_ad13_b446_d0eb_abe4_1f88_556f;

        #200;
        key = 128'h7d3d_4e3a_1c2b_0e0c_4d32_42d9_0e26_61f8;
        state = 128'hf210_0592_1fa9_9300_1924_487e_0f3c_35df;

        #200;
        key = 128'hefd1_3492_9160_737e_fb47_29c6_8c05_f5ff;
        state = 128'hd3cb_0a30_a1fb_d5a7_e33c_2606_9e24_edfb;

        #200;
        key = 128'he64a_14b2_c0c3_d244_aac3_03b0_3e58_e8f0;
        state = 128'hcf4f_c53b_bda7_df17_e291_553d_16e6_daa2;

        #200;
        key = 128'h5383_f82b_b0e3_b01f_3a10_d37c_0316_7cd8;
        state = 128'ha8c5_6d4b_b67b_b144_7e7d_c4f6_7d7c_7d59;

        #200;
        key = 128'hf9b6_4930_9b46_d4fe_3beb_f43f_cb2a_35f2;
        state = 128'hbf6a_b11d_7fd8_3d02_183f_e76a_6222_f1ed;

        #200;
        key = 128'h3860_2096_ec22_4a97_3530_6608_94a7_6d75;
        state = 128'h7855_a46a_a6f0_8ee7_de81_f2f1_a9d1_d814;

        #200;
        key = 128'h465f_cc4c_4b33_7fdb_3a80_5bb6_3f2c_a21c;
        state = 128'hdcb2_cfc5_930f_53f9_26b4_922b_45b4_7c97;

        #200;
        key = 128'h2b36_4603_ffab_f89d_19d8_5e34_a1f8_322d;
        state = 128'h9e9d_8c75_43c9_160e_252b_5dae_6385_0a33;

        #200;
        key = 128'h5766_11e7_f3b1_8bfb_2744_61b2_0de7_4cd9;
        state = 128'h16da_4fe2_6d8b_66bb_5872_56d1_348d_da4d;

        #200;
        key = 128'hf45e_6557_bcc5_3f89_2924_5c28_52d6_a81b;
        state = 128'h59c1_6d3d_9140_17a8_472f_2ee7_a10c_356d;

        #200;
        key = 128'ha278_b09c_6c77_e1bf_2e3a_eff2_b178_b9bf;
        state = 128'h9e54_fc09_dd26_0cfb_cb07_8251_b9e0_0a23;

        #200;
        key = 128'h4e9a_f3f4_61ab_c9f2_4fe5_afd6_fc9e_b955;
        state = 128'h1193_8d67_c683_5f37_a214_c491_3c82_62bc;

        #200;
        key = 128'h6746_4467_f073_a18f_3999_2f89_ce20_79f3;
        state = 128'h149d_a85e_8809_1c2b_4c8e_9b43_a9c0_830c;

        #200;
        key = 128'h14be_cad5_d196_475e_3aa4_e88e_0511_ce64;
        state = 128'h2c25_5e04_b5e4_20b3_77e1_6562_4bec_3ad4;

        #200;
        key = 128'h556e_278f_3ea7_a936_d4c3_13b6_4a41_979f;
        state = 128'h0c6d_7205_ee2c_c26a_de76_98eb_694b_3d57;

        #200;
        key = 128'hec39_03d3_b102_34cb_b437_e67e_613a_2070;
        state = 128'h0e90_6d80_f5b8_9c52_c618_6ecb_5f47_89a9;

        #200;
        key = 128'h094b_7497_bd19_f502_8ecb_0cfc_488e_1663;
        state = 128'h2735_3af8_281f_9528_1c04_1bc4_569d_8380;

        #200;
        key = 128'h3dc8_57bd_bff9_2450_3b79_2cca_5c9a_acbf;
        state = 128'h2743_c021_2b68_9a2c_59b6_c6d8_6053_d223;

        #200;
        key = 128'h9861_e296_e8de_7005_1584_cd1c_18eb_6f43;
        state = 128'hc785_2e72_ad99_c72c_6dcd_9ca4_92db_8a67;

        #200;
        key = 128'h03fd_71d6_65ec_c1a8_5e4b_d6ab_85ae_4f8a;
        state = 128'h1358_0623_72a3_f225_5977_0d82_b9d5_0476;

        #200;
        key = 128'h496a_c438_0223_cb86_035c_7b49_6341_88a9;
        state = 128'h2757_98d3_bf95_af56_7d8e_bb60_2d67_f435;

        #200;
        key = 128'ha00e_42b3_15b7_5648_93ba_147a_496e_215a;
        state = 128'hea33_1ff9_b7cf_d074_9748_d459_50de_b2f9;

        #200;
        key = 128'h9139_6505_90bd_157d_dc16_897b_354f_844d;
        state = 128'hfd51_0fbf_fb01_f5fa_7885_5744_2037_4e93;

        #200;
        key = 128'h6437_2e6c_6a30_4bbb_9c83_eafe_f445_5e3e;
        state = 128'ha336_dccf_a759_d4ae_edc4_4556_3f2e_a3d9;

        #200;
        key = 128'h472a_be1a_2b09_b3a7_63ad_b2d2_bb57_1f44;
        state = 128'hed7e_4247_3a87_f4c9_9bcc_7e1c_cc68_7469;

        #200;
        key = 128'h47b7_1b8a_41c0_ad92_51cc_6397_ea71_dc16;
        state = 128'hc99f_ecf6_b5d1_4bbd_89e6_fec8_b971_fa68;

        #200;
        key = 128'ha5a1_5acc_e1b9_bc3c_5f46_e7cb_61a8_ec1e;
        state = 128'h2523_e86f_9ac0_a3ad_5bda_fbc1_537b_8e04;

        #200;
        key = 128'haa10_ea8e_b075_ce23_f22f_c27b_74dc_8d47;
        state = 128'h964d_4a37_4010_e79b_848b_5b69_e6c9_eab9;

        #200;
        key = 128'h6325_ce44_0921_a29d_038b_bc29_342d_f208;
        state = 128'h1013_1d20_ae00_2865_50d5_23e7_4dd1_937b;

        #200;
        key = 128'h20e6_a136_73ae_5805_b90e_23c2_d2d0_7d62;
        state = 128'h4883_caa5_81b6_08ba_d6ad_1bae_fe3d_0c28;

        #200;
        key = 128'ha104_3219_e6dd_88f4_ebff_fd8d_d3b2_7e24;
        state = 128'h6d4f_2bf1_047f_f56d_ad0b_e342_b978_6075;

        #200;
        key = 128'hab51_77b0_522c_6f71_8e56_5dff_c5b6_5af5;
        state = 128'haff5_781f_ced5_abd1_9543_d96d_38a6_2f4f;

        #200;
        key = 128'h7387_d34f_0813_00d6_5181_fbcd_0c17_32e6;
        state = 128'ha7e5_d094_0ad8_d951_7521_0876_8537_98fd;

        #200;
        key = 128'h42c4_48d4_080c_fc75_1c47_ba14_e9be_b6f3;
        state = 128'h9737_1f62_9cdd_3380_fa28_33de_dfd1_a22e;

        #200;
        key = 128'h685d_2f51_5674_d0e3_ffde_ec21_1462_7ea8;
        state = 128'h9314_08b2_c26a_e1d2_0344_7f57_2c35_5b4e;

        #200;
        key = 128'h20a0_d5d1_74d7_6987_edb5_8160_4203_1e42;
        state = 128'hf6b7_1c36_3e77_62c0_156d_61e1_d60c_50a2;

        #200;
        key = 128'hf5a3_fae8_b702_0774_ed2a_ea9e_b410_c2a1;
        state = 128'h866d_0ea2_dfb1_ef3e_20ba_3a5e_5873_4c17;

        #200;
        key = 128'h5ace_393f_6950_b761_b5dc_e546_9555_9dc0;
        state = 128'hbde1_4689_7dc5_b21b_7464_775a_e3e0_0089;

        #200;
        key = 128'h4004_510a_998e_ec12_0477_efba_ead1_d6af;
        state = 128'ha95d_3f46_1cd8_8fb2_b0e1_6799_da9d_2e50;

        #200;
        key = 128'h9d12_69fa_826a_79f4_a1fc_cacc_ec2f_3943;
        state = 128'h7e2e_c754_a391_1f9a_bb9c_df1a_4264_7927;

        #200;
        key = 128'hca98_3699_cb79_7e0e_90cf_8b9e_971f_67ad;
        state = 128'h97bd_d625_eefe_aeaf_2707_4efa_1fa8_7f21;

        #200;
        key = 128'h6a05_a050_a483_431d_55b6_76bd_3ab8_bfcc;
        state = 128'ha0de_74e6_b23c_84d0_22f5_0b0f_c6ee_3e57;

        #200;
        key = 128'hb606_866e_a972_cba3_b4bf_ee80_8b47_1566;
        state = 128'h1aa8_640e_46da_d6c1_c931_d018_b039_a07c;

        #200;
        key = 128'h12e5_a2a3_9761_f82b_b391_5006_1edd_9cd2;
        state = 128'h0ee1_ed15_626d_0d74_0844_22c8_8c77_6050;

        #200;
        key = 128'h5b32_8c3a_ca6a_ebb0_aa17_0a8a_524e_b73f;
        state = 128'h8b2a_db03_3685_7f74_d3b2_0ff8_fbc0_171d;

        #200;
        key = 128'h4aad_0727_f819_5968_8109_a17c_9eb3_5566;
        state = 128'h5729_2af2_53c4_75c9_68c5_c74e_fba7_0b05;

        #200;
        key = 128'h8fde_5efd_ed4a_c2d8_b070_0f1f_08f2_4b1b;
        state = 128'h9243_798c_3674_eb11_4b5f_20a5_3cc4_111e;

        #200;
        key = 128'hef8b_6dde_1c1b_cc2f_8a33_9abf_0701_d7ca;
        state = 128'h82ac_fc9e_bcdc_81a2_f322_1376_2def_d101;

        #200;
        key = 128'ha449_c782_2b89_7fb7_6b95_a2b8_3947_6a25;
        state = 128'hd086_fa0a_86e5_915e_8306_e681_4b2a_5714;

        #200;
        key = 128'hab0f_7982_0272_864a_c143_d434_2fd1_4815;
        state = 128'heca2_11e6_97b4_6739_54ff_cd19_b6b9_e16d;

        #200;
        key = 128'h42da_fa3c_7d1d_c108_869e_7690_de81_2960;
        state = 128'h1503_2406_adaa_b3c1_b9c1_1f40_d432_12c0;

        #200;
        key = 128'h0b1b_805d_bf35_a5a8_0a72_97c5_1b3b_b718;
        state = 128'h295f_94d1_6e48_6fee_6bf2_a4b9_37d9_33ab;

        #200;
        key = 128'h5160_c685_ce4d_7ca3_5884_8580_ea15_fcce;
        state = 128'h1cda_8aa4_3e52_8450_3161_5df5_9719_0f87;

        #200;
        key = 128'h56a9_1bbf_4d5a_5830_d90e_a6b9_5810_8589;
        state = 128'h6199_8aa7_a013_7796_bd80_5519_11b5_0d4b;

        #200;
        key = 128'hd717_9d46_e60c_5613_db9c_77cf_7324_13b6;
        state = 128'h65f1_e4ee_4791_46f3_dc35_66a8_e0c4_04db;

        #200;
        key = 128'hb30f_b4f8_abcf_900d_dad4_d914_e105_4ef1;
        state = 128'hf98e_e872_9d38_59cf_3bc5_2d0e_fd05_954e;

        #200;
        key = 128'h946f_7513_8065_501e_6428_3296_0852_a460;
        state = 128'hb928_d4ff_86d4_acc5_ba4c_2cea_6ae5_f1d2;

        #200;
        key = 128'h4572_67b8_16cb_3b0a_33f1_a44a_1f01_047a;
        state = 128'h8ac5_c6b0_8155_2f74_b16d_dfa1_9c48_e81f;

        #200;
        key = 128'h09d4_21f7_2dbb_6fbc_b1da_8fc8_adfa_998c;
        state = 128'h4cf0_c7c2_1076_05e5_84bc_8eb7_2d30_f4b9;

        #200;
        key = 128'h3284_cfe7_6b4e_60c2_89f1_84f7_ea89_b35a;
        state = 128'hce13_5476_9f7e_824b_885f_821c_abf5_1c35;

        #200;
        key = 128'hcc5a_0475_c773_87b2_c926_059b_b3c4_e30e;
        state = 128'hcb86_4218_3cdf_c97f_9d2f_4ef7_59f4_1ba1;

        #200;
        key = 128'h37a6_6a35_58ac_028f_8205_3b8b_ed0d_21c9;
        state = 128'ha3c6_74a4_0c1d_a4cc_e621_837c_9b72_3bce;

        #200;
        key = 128'h5895_e68a_8367_ed6a_9607_24f7_ea80_8351;
        state = 128'hb3a9_7bbf_448c_9715_619b_f518_1ec5_f4a3;

        #200;
        key = 128'h6418_9df6_e598_f7dd_9c5a_ef9d_5611_ef4a;
        state = 128'hface_143b_84c1_f4c9_d3dd_f3a5_877b_a521;

        #200;
        key = 128'h2a89_3b1f_538b_14c1_c501_304d_6f00_c144;
        state = 128'hf2ff_5dd7_edb9_6163_6b33_c413_e5cd_1196;

        #200;
        key = 128'h8a6b_0dee_44cb_c30b_ed46_bbbc_47c8_35df;
        state = 128'h55f5_6c9d_c875_7cdd_47bb_e61b_a3a7_16b9;

        #200;
        key = 128'h66a3_d968_0282_9cfa_e237_8888_0714_e2c4;
        state = 128'hd7e2_6b9a_b8f6_2e20_3f32_485e_c554_384a;

        #200;
        key = 128'haeae_a269_72b7_bdaa_8ab1_6a91_be4a_c816;
        state = 128'h1dde_6de9_68b6_3aae_29d2_e3e0_2cf6_0542;

        #200;
        key = 128'h1411_ee68_464a_d221_2037_0c0a_45b3_f36a;
        state = 128'hf2da_bb67_3c6f_68f3_ca8e_b343_e85c_6624;

        #200;
        key = 128'h2d45_81d0_bc4c_bd79_742c_6cd5_321a_0796;
        state = 128'h4b6d_f77b_0ab6_1fa7_4c22_63e3_09fc_ce3c;

        #200;
        key = 128'h4ac7_7aaa_992a_1b26_911f_9ade_e7a3_b8e4;
        state = 128'h8519_4a3c_f914_f8ae_47af_8982_d2bf_8bf0;

        #200;
        key = 128'h7080_870a_0851_980a_444e_e0d7_bed8_2cd6;
        state = 128'h2768_e254_f2d2_3828_e500_7392_1c1e_1ce8;

        #200;
        key = 128'he94e_ada2_98b7_a9bb_fb62_2978_2a71_cb99;
        state = 128'h3c77_c94e_f8b4_ebbb_6df2_6ee9_0504_a3d0;

        #200;
        key = 128'hdf84_5054_8d81_79a2_f1fd_bbe1_7c79_1777;
        state = 128'h71ef_a414_cade_95c6_8677_dd74_d082_3462;

        #200;
        key = 128'h123f_c89b_2da7_a6ca_01af_c9c7_09e9_b29c;
        state = 128'h4981_38eb_10fa_ff1d_33e9_013b_09c1_35e6;

        #200;
        key = 128'hd142_11aa_c6f4_506c_7ec2_e396_b8dc_dca2;
        state = 128'hebc0_bf75_77a8_fdb2_77c4_2be7_c898_5238;

        #200;
        key = 128'h39a6_360b_661a_e26d_ba7c_7802_f80a_f01c;
        state = 128'h2e7a_cdcd_48bc_a9bf_2d11_51ce_a38f_4200;

        #200;
        key = 128'h3e86_f527_4a1e_4c14_f4e0_8a8e_83f5_f494;
        state = 128'h96b8_17f0_840a_dd63_8618_0bbd_f467_a00d;

        #200;
        key = 128'h7fb2_5197_d7ce_c6d2_cc65_c488_9571_7c35;
        state = 128'h9a2a_fe15_5105_0252_f312_44f6_faf8_2fc0;

        #200;
        key = 128'haebc_803a_1e94_1df1_c37f_65eb_d900_2d5c;
        state = 128'h367f_d3fd_353e_edd1_4245_f836_b9d4_7d97;

        #200;
        key = 128'h418e_ec35_d58e_88bf_bff7_4f20_8aa7_3dd5;
        state = 128'h8bbb_9504_b3a4_8de5_0ea6_d9ac_b11a_83c7;

        #200;
        key = 128'ha867_dd43_cdfc_01b6_95ae_b63e_43f7_0839;
        state = 128'hf578_dc29_8652_2d0d_bf63_2532_7467_035e;

        #200;
        key = 128'h69a9_c768_b3fa_dcab_8098_61b7_0816_8c1f;
        state = 128'hb476_2b60_3111_80fb_74b6_6407_d4de_6ce9;

        #200;
        key = 128'h4ac4_db99_41c2_22de_7891_62b5_ca66_38ed;
        state = 128'hf634_c222_8009_c4d1_d134_cbca_539a_b774;

        #200;
        key = 128'h140f_63cd_de5f_c923_ba40_dc1f_e823_c2aa;
        state = 128'h7f2d_11ff_077c_0ab1_00da_dd09_6af5_fca5;

        #200;
        key = 128'h29ab_4f2a_3cf4_1299_63cd_8810_e414_d8a6;
        state = 128'heed6_bd7c_9ae7_2afd_9d83_b366_aa33_1b3d;

        #200;
        key = 128'h5742_04e3_86ad_a220_e0bb_09ff_479e_7ee1;
        state = 128'h8bb3_e572_48df_8437_3028_6cd0_fb31_8ec0;

        #200;
        key = 128'h6299_353a_3559_cd6b_4a46_a33a_36d4_3a51;
        state = 128'hafd3_6ea6_3729_5d43_c2d8_33dd_8b9b_10a2;

        #200;
        key = 128'hbf6f_b886_3183_b6a6_f4bd_6007_ff60_6e8c;
        state = 128'h4d19_2a3f_c480_24b6_a91b_91ca_96be_b65c;

        #200;
        key = 128'h2b1c_aa0a_2fad_c1e5_733a_337c_ef3c_b9cc;
        state = 128'h8e32_889c_a94d_b841_df48_e8f5_a016_6039;

        #200;
        key = 128'h9c97_c67e_555c_70e2_3290_2d2d_302f_3ea5;
        state = 128'h9bbc_3568_48c5_dccf_b3cc_445b_a2ac_11b1;

        #200;
        key = 128'hb06b_a0e8_de4f_50d2_33d5_66f1_6ff8_bee9;
        state = 128'hd02b_f069_7a8f_44cd_067f_4183_af04_a084;

        #200;
        key = 128'h3995_af23_2240_29de_06d6_42ca_25f2_b6d0;
        state = 128'hf976_8e15_dfbe_1396_ca26_9cf3_de5e_81ae;

        #200;
        key = 128'h5e7b_5bf3_8e63_fbb2_6918_6e85_010f_3562;
        state = 128'h628e_41c6_4f34_94b2_6f5c_17a1_3003_3392;

        #200;
        key = 128'h2a56_929b_85ca_31ad_4e0c_405f_55bc_116e;
        state = 128'hef2e_3260_1410_c9c0_7e1c_251e_a519_b825;

        #200;
        key = 128'hce1c_8877_473e_197f_496b_f810_48dd_8e7f;
        state = 128'hf5d9_00af_85b4_b51d_2d71_7772_2b2c_cbad;

        #200;
        key = 128'hc84b_3f61_f9f1_b688_27e0_bc43_6b6a_b9f5;
        state = 128'h9708_a25e_2e96_b90c_52a2_5108_7905_20eb;

        #200;
        key = 128'h0f78_f206_9ce7_92fa_69ba_440d_48e5_a152;
        state = 128'hf934_1ff0_dbb5_c745_97ba_1eb0_a103_4a75;

        #200;
        key = 128'hafe7_3d64_529b_7248_accb_47ef_cea5_3de7;
        state = 128'h952d_d715_058f_4854_4b28_fbfd_b363_006a;

        #200;
        key = 128'h0f95_2344_6cb3_2071_2af4_c31a_a2fc_aa48;
        state = 128'hb25d_2853_b321_f34e_df2a_bb63_8de9_44d1;

        #200;
        key = 128'h892f_1057_9a0c_36a5_8130_368b_61e5_f5a5;
        state = 128'h97ea_2ec8_db54_1468_2b7f_f12e_c345_8aeb;

        #200;
        key = 128'ha47c_af77_8faa_2f30_0dc2_e065_c0d4_81b8;
        state = 128'hbfbc_101a_0e3c_c390_f1eb_3895_d6cc_9c38;

        #200;
        key = 128'h2a0f_320c_3ca3_90f8_43a6_0252_7347_eaf0;
        state = 128'h70fa_a636_4807_cb38_d470_16b9_c62c_7a57;

        #200;
        key = 128'h4009_ee1a_f8d2_3809_6c59_55e6_ff6d_66a3;
        state = 128'h1ca0_ea4f_acfa_52ea_4830_d163_98c0_9959;

        #200;
        key = 128'h1266_e3ba_7daf_342e_3879_b3d4_6282_2a4f;
        state = 128'h2fe6_e38d_430a_34e9_0e10_1ac5_c57c_cbff;

        #200;
        key = 128'h1211_0d1e_272b_a555_af78_0476_5d53_7c2e;
        state = 128'hb098_f198_fb62_9360_a6b6_3241_c06b_c50e;

        #200;
        key = 128'h9ba1_6db2_90cd_83cd_b36b_f38d_643e_9221;
        state = 128'h2199_b0b2_90db_a752_9b28_1e15_901a_b172;

        #200;
        key = 128'h7a14_b972_8ffa_89e6_1318_d98d_0a0f_3b16;
        state = 128'h9860_4199_75a8_ec18_e3d2_95b5_bbf2_a8f6;

        #200;
        key = 128'hd85c_0b31_20ec_0499_6287_cc85_9a39_bb0c;
        state = 128'h8a77_44fe_94d8_53dc_d288_7cd8_c89d_9b30;

        #200;
        key = 128'hdab2_bab2_aa1c_cdfb_17d5_b7ce_2824_88fa;
        state = 128'hd1b2_851d_63de_fa2c_2e58_57e7_a3c7_098f;

        #200;
        key = 128'h4ce6_9973_4a8d_2f7c_b90d_57ea_8328_e6b7;
        state = 128'h5dc7_762d_ca7d_6912_6fa4_13e8_fe4d_e00c;

        #200;
        key = 128'h481e_1286_f6c9_0ecc_b0d5_c3e9_e7ff_725b;
        state = 128'h59a2_dcbc_fd04_0261_b940_1c69_02c9_99f8;

        #200;
        key = 128'he469_efe9_bf02_c95f_929b_b399_1841_873d;
        state = 128'h8de2_94fa_2297_81bd_08c1_0b36_508d_56c0;

        #200;
        key = 128'ha5a6_2179_3021_f54b_8676_1c8d_e292_a6af;
        state = 128'h49d5_d82d_14b7_8108_394b_9e76_9a5a_8219;

        #200;
        key = 128'h2ede_519b_ffc3_6575_0d60_a461_0894_81ca;
        state = 128'h4d10_5e67_9e57_65b8_18a8_a7a4_944d_d20b;

        #200;
        key = 128'h35fb_0fcf_20e2_7ee9_0588_4b27_411a_38c8;
        state = 128'h9438_9207_c7d8_d97d_24bd_f8bd_6b18_ea8f;

        #200;
        key = 128'hd028_bc8c_9d58_e4aa_6374_4d17_b774_7977;
        state = 128'hef10_a087_8caa_3fa7_e55a_e44c_896f_883f;

        #200;
        key = 128'hb224_9f96_6959_bf02_e85f_77f9_8b3c_a8c2;
        state = 128'h3c3a_8096_f407_0f87_3157_10f8_8f1c_8c2b;

        #200;
        key = 128'hf0d9_c1e8_7e2d_8449_c3c2_a149_43ee_1567;
        state = 128'h60bf_a49f_a221_eb7d_03c5_8df7_b9bc_e8df;

        #200;
        key = 128'hf782_fdad_7883_765d_32de_9e70_fd8e_9667;
        state = 128'hbfce_3fdf_2f19_31df_4769_1986_9658_fdb5;

        #200;
        key = 128'had16_5d5c_c9fe_39f2_417e_9c5b_ac5f_9659;
        state = 128'h44c3_546b_e8c0_717c_abf4_fd77_5b56_0683;

        #200;
        key = 128'hce76_051b_2ee6_6797_34e2_0459_0d3d_61c1;
        state = 128'h324b_b2fb_184a_74a0_3c3b_5d89_0050_a3db;

        #200;
        key = 128'h2983_ec15_cc80_4a32_94bf_c9da_3bce_6914;
        state = 128'h2734_c99d_1291_1496_98f9_367d_f0a2_1ec9;

        #200;
        key = 128'h004b_eb37_458d_7db1_3130_5ad3_efde_b1f3;
        state = 128'h1760_2962_76bc_492f_8471_7207_0314_ae24;

        #200;
        key = 128'hd03d_41e7_3058_30fb_a9d8_edfc_2bd7_493a;
        state = 128'hd1c5_4af0_1883_37bc_ad7d_8e71_6eb2_ac34;

        #200;
        key = 128'hd040_a1b8_f3a7_31e9_2bad_6dac_c637_12df;
        state = 128'ha053_50f8_06cc_d913_32e6_777c_060f_f94e;

        #200;
        key = 128'h393f_2049_070e_eb70_e492_b6b3_26f7_ccc1;
        state = 128'h7dc8_45e9_036c_66da_dea4_49df_57e4_a505;

        #200;
        key = 128'h3d4e_a955_e1a0_68c7_f717_0800_e204_9752;
        state = 128'h8ab9_278b_b2b9_13a8_4a04_f20f_8218_819c;

        #200;
        key = 128'h90c3_1851_7c5a_6aff_ebd8_3cb0_1f20_99ae;
        state = 128'h8d07_96e3_e61b_c49e_0ddd_db83_2bba_6d16;

        #200;
        key = 128'hdaa2_6df4_492b_27d3_425a_c1d5_8980_55f8;
        state = 128'h4484_bbf8_7a2e_76ae_c88a_047b_d3b7_5460;

        #200;
        key = 128'h8d90_dadb_c040_78fe_ad6b_8e43_79fc_58e2;
        state = 128'h0ce8_d124_ce26_e775_2951_c90d_d659_5dd3;

        #200;
        key = 128'h49f5_db7f_db27_be34_7b9c_423c_257a_7b4b;
        state = 128'h734d_881d_f5e4_b1d3_4909_4feb_9995_6cb9;

        #200;
        key = 128'ha607_3ff6_8609_b4c0_e7fc_d3c9_96ce_715e;
        state = 128'h499e_bf14_6649_57d8_44ef_a8e0_1d96_b04f;

        #200;
        key = 128'heef5_c1a5_fbde_22ad_9be0_123d_bde5_3dd8;
        state = 128'h5975_1549_77ae_009e_66a7_b54a_d574_4854;

        #200;
        key = 128'hb0f2_75fa_96ab_72d7_35ec_01e2_b94a_8dcb;
        state = 128'h5d63_d82d_19b2_20e2_da53_280f_1512_5c14;

        #200;
        key = 128'h004e_8843_edb6_7260_855f_bba3_3c13_af02;
        state = 128'h87c0_fb85_6034_c1c2_1845_e7f3_72a1_076b;

        #200;
        key = 128'hca97_2e71_1a7d_73e2_0ed6_c46d_7325_10bc;
        state = 128'h8afe_6be8_60e6_6e25_4621_7776_e1cb_7278;

        #200;
        key = 128'h9b80_8dc7_7dad_d773_5d73_d01e_17c8_332b;
        state = 128'h0341_5493_973b_1d03_1719_f5b4_d385_9504;

        #200;
        key = 128'haa98_614d_8d73_7229_15ab_5adb_cf7a_9a4c;
        state = 128'h190d_44b9_7386_7b6e_6252_4a40_f4d0_44b3;

        #200;
        key = 128'hb3b5_4ed4_cc0a_59f1_2a04_dd26_dd37_f7f4;
        state = 128'h5f04_b306_49f6_ffe0_c497_1b83_ab1b_3d60;

        #200;
        key = 128'h7d09_ee0f_a7dc_3c4b_a2cd_bc22_4be8_ff10;
        state = 128'hd611_26c6_c273_624c_1fe7_4256_ffb3_60a7;

        #200;
        key = 128'hd004_73c1_2698_8a7c_65ab_3bee_da0c_8d23;
        state = 128'hae01_83ef_7073_46f1_eda9_9901_9233_ece8;

        #200;
        key = 128'h6087_1a8e_da55_2c8e_b24e_d701_1c3e_a996;
        state = 128'h0066_b230_a37a_b573_b5dc_7068_b0f3_bf4b;

        #200;
        key = 128'h9d43_e92c_a05c_f76e_648d_18af_6c29_5aac;
        state = 128'h323b_7ac6_3274_f43a_af07_404e_9e97_c1ad;

        #200;
        key = 128'h4d0f_5a5f_64b1_ef7c_caba_cd37_fb72_1a17;
        state = 128'h581c_1f07_c8d4_f828_b50a_fe93_9998_4269;

        #200;
        key = 128'hdad8_b7ed_3264_95b0_d4d8_2997_eb06_1eae;
        state = 128'hc775_f1a9_55c6_3de7_dc14_40f7_0a25_6c0e;

        #200;
        key = 128'hf65e_d498_464a_8579_29f0_3fc1_aef3_3ac2;
        state = 128'h03ab_d2ff_17f6_aa2c_961a_32e0_6323_047b;

        #200;
        key = 128'ha1c2_1448_a737_86ee_d106_bf3b_643b_df54;
        state = 128'h8ac2_826f_8509_49cf_c1c7_7821_b3c0_1329;

        #200;
        key = 128'hf78e_28df_0e7b_814f_c5b4_bb0f_95c1_5257;
        state = 128'h8109_3c82_fd94_9c6f_e94f_4f64_ebbc_a567;

        #200;
        key = 128'h249a_0019_d6dd_d060_315a_1b4b_e693_10d4;
        state = 128'h6b8a_7985_1cf3_8016_b368_6675_b11b_7ef5;

        #200;
        key = 128'habf4_55a0_18fa_f514_fda7_a6ae_a084_cd72;
        state = 128'h550c_66c4_5bb0_0dbf_c383_0b49_c463_d510;

        #200;
        key = 128'h662f_892f_a80d_3ee6_a2f8_b2d3_b84e_704b;
        state = 128'h38ba_0fe6_a763_85d9_3270_b666_1a49_5079;

        #200;
        key = 128'h8dc6_4862_5ab2_e45f_04fc_bd46_8129_2ba8;
        state = 128'h93a0_a8aa_2415_e6ca_520e_ed09_82b3_e31e;

        #200;
        key = 128'hee6c_c0c1_4197_cd09_1dc3_c4c2_d53f_1968;
        state = 128'hfd13_ccef_bff5_aa07_59ed_0ae7_bb26_333b;

        #200;
        key = 128'ha613_3503_2df0_641e_b52d_f69e_aa8b_53c5;
        state = 128'hf65a_413e_e4f0_ad1c_5da6_2a36_ac3c_bca3;

        #200;
        key = 128'h9c38_c982_2581_0dcf_f756_a286_0b1c_bc20;
        state = 128'ha00c_872e_3006_03c1_5642_f28a_c9d5_f392;

        #200;
        key = 128'hcae4_4821_35f5_824e_91d2_624e_3d6c_c78f;
        state = 128'hb87c_5b5d_0e3c_c704_db36_9a11_1cef_1832;

        #200;
        key = 128'h467e_238b_a594_4509_64ff_f124_c23b_0510;
        state = 128'h0f9a_a989_09d3_9d09_c61e_84a9_9465_323e;

        #200;
        key = 128'hc81a_3846_f3b8_3a73_0281_1efe_7a13_a952;
        state = 128'h68d2_e545_52f1_2539_86b8_5ee5_7327_c1ce;

        #200;
        key = 128'h2f15_2702_6b77_2bec_bb26_7c97_dcdf_6219;
        state = 128'h412f_ffb6_33e8_414d_c189_d39f_3431_0f02;

        #200;
        key = 128'h13c4_638b_7fb2_9a29_540a_4e7c_94f1_bf9c;
        state = 128'hfabe_0bae_5c02_127d_361c_daf0_1ae0_f994;

        #200;
        key = 128'h6b58_387c_1b6b_74ab_a033_63fc_d5e7_87b1;
        state = 128'h5c49_47e8_7abc_8d78_b0b7_6c15_22e1_5b65;

        #200;
        key = 128'hcd8c_edc5_8c39_21c0_5b29_822a_eb02_34b2;
        state = 128'hc42c_c6d3_e328_38f9_503c_3f29_046a_e3fd;

        #200;
        key = 128'h2433_1913_6eaf_eeb2_da79_c97d_06db_f04c;
        state = 128'h28d7_241a_1e3f_22bb_03df_5dcb_68c1_708d;

        #200;
        key = 128'ha61a_1abd_b378_725b_affa_1a24_ebec_f0b5;
        state = 128'hc13d_dc39_3786_ecae_358d_6291_7bf7_76e3;

        #200;
        key = 128'ha7b9_cbbd_037d_78a5_cb66_311a_65ef_38b1;
        state = 128'h3c18_98d2_aaa6_4b65_a35a_a4f1_142b_fe51;

        #200;
        key = 128'hd612_7f98_12b9_9c29_286f_e91a_f28f_52c3;
        state = 128'h55fc_0f0f_ee83_ac36_b475_26b6_2b51_6478;

        #200;
        key = 128'h08f4_31ec_3bd7_04e8_fe99_a416_9bc4_1b78;
        state = 128'hf7df_82e9_2331_0754_c9f9_5509_c9ca_4374;

        #200;
        key = 128'he7f8_55f3_b3b5_a515_794d_4be2_b6f2_6c91;
        state = 128'h51ee_e5fb_9de6_fbe9_992f_8f3d_b98e_dc81;

        #200;
        key = 128'h0638_1366_f3c4_30c9_44c2_012e_3992_2b93;
        state = 128'h6fdf_5310_998b_ec85_4c32_d2fe_482e_3b3e;

        #200;
        key = 128'hd32b_ddc3_af37_ec95_e5b4_0b9e_0cce_1e1b;
        state = 128'h9bbf_6424_1893_ae6f_bace_112d_51f8_df12;

        #200;
        key = 128'hcc76_9e18_cc7d_55a9_0e25_8019_46f2_108e;
        state = 128'hc632_e523_f9e3_9c19_e471_dec0_5157_eda4;

        #200;
        key = 128'h8146_d205_2271_2ad7_adc7_8000_7ba6_0216;
        state = 128'h73cc_d2cf_01c8_0a8d_4eda_a8c9_1911_726b;

        #200;
        key = 128'h3cc4_ead5_798d_4c2e_6dea_00ab_8c6f_69d5;
        state = 128'he8af_4ceb_0ee9_3019_7b5c_6060_e7d8_6679;

        #200;
        key = 128'h541d_13de_4895_9e0a_60e3_2c91_d000_76ae;
        state = 128'ha341_d1ed_fa89_381d_b7b6_1c44_1065_c1eb;

        #200;
        key = 128'h2348_affb_64f7_19fd_3c02_95d0_e391_11c9;
        state = 128'h33fb_a152_1018_2f4e_8ce2_8dee_26ef_0ec0;

        #200;
        key = 128'h691a_c063_9327_d89f_14d5_c178_4b93_b3e5;
        state = 128'hdbb2_2566_39df_de17_54b8_4be8_2d5a_f7c3;

        #200;
        key = 128'hb73f_f506_9ff2_9102_63cb_a23b_ddb0_7777;
        state = 128'h947d_c63d_7094_ccbb_226c_0298_17c1_e4ea;

        #200;
        key = 128'h00ce_3058_cd84_1eac_1051_c0ba_0d40_f344;
        state = 128'h1b6e_0890_64c4_7398_b1c4_9486_a285_1974;

        #200;
        key = 128'hfd68_a520_16c7_e2d4_454f_3ffb_63fa_fb44;
        state = 128'hb399_3871_7dcb_8ec8_6085_5871_4875_f180;

        #200;
        key = 128'h3319_ce3e_9e41_681e_dddc_456f_f2a1_d8eb;
        state = 128'heec1_0606_7dd8_331c_7ac0_2e3f_17ea_e2ce;

        #200;
        key = 128'h5d3f_0f54_b49e_29f4_c02c_6606_40c8_6299;
        state = 128'h8c11_0f0a_db0b_1702_9f29_9266_f341_5e0a;

        #200;
        key = 128'hc906_fe0e_aa29_977b_1e58_cf9d_6187_1f51;
        state = 128'h7c6c_9d3e_a6d8_a279_0d4c_238a_677f_c63a;

        #200;
        key = 128'h4fa9_7216_9e56_65ff_a37b_98ea_512d_bdae;
        state = 128'h7c5b_c17e_31d4_9cab_c4ef_ff04_eeec_f35d;

        #200;
        key = 128'h0d02_67c5_05a6_a6de_d17c_9497_3c0f_ec2d;
        state = 128'h4512_8a3a_28bb_2b69_65b3_05c9_b404_c77b;

        #200;
        key = 128'h39d5_fb52_23ac_e7f0_6ae6_f265_1a1d_e811;
        state = 128'h329f_51c6_8d81_34a0_bc56_b539_e098_34ca;

        #200;
        key = 128'hb63b_3020_de18_5354_8af8_4f34_397a_3243;
        state = 128'h5ea9_6753_b2f8_7032_76db_3672_716f_8113;

        #200;
        key = 128'h8445_38ee_2696_fa62_1473_d47b_4e07_8fee;
        state = 128'h4009_7a1a_be48_3409_6f7c_e763_2ac4_0870;

        #200;
        key = 128'ha938_e820_0ba3_435f_da8c_9d26_901a_e2db;
        state = 128'h2bf8_b232_2ee9_5417_79e2_0468_028d_887e;

        #200;
        key = 128'hcaaf_4f8e_5821_6030_06e7_d28c_3522_2c14;
        state = 128'hc83f_8aa4_3098_d17a_3982_6ea2_a2dc_4ab7;

        #200;
        key = 128'h9e87_abaf_02a0_259c_f13f_044d_584c_9f82;
        state = 128'h89cc_ddf9_8d4e_46c6_7946_41b3_c165_fe39;

        #200;
        key = 128'h2930_3f61_e429_1936_a11c_adf6_340c_804a;
        state = 128'h19db_c873_ccf7_4ae7_7011_bd65_7e2b_51a8;

        #200;
        key = 128'h7771_0fa8_f731_f55f_b894_9600_32ca_efca;
        state = 128'hc485_687b_f214_0a2d_4caf_e7b3_2bb1_dd2b;

        #200;
        key = 128'hcfc4_0b81_449f_c241_c57f_f43f_e4ed_8511;
        state = 128'h7980_2627_5a5e_a498_d45b_a59b_4a10_43fa;

        #200;
        key = 128'hf623_65cc_de9b_df4c_35de_38ae_5111_3684;
        state = 128'hb387_698e_0c1d_3367_fc82_2033_6832_129f;

        #200;
        key = 128'h7627_217a_c132_60db_2142_3b94_3753_931f;
        state = 128'h5322_f804_4833_f8f4_09af_a961_6819_2364;

        #200;
        key = 128'h93d4_5588_597e_611f_2500_cfbd_0910_2344;
        state = 128'hf75b_4bc4_221b_02bc_bfd5_78de_7af5_39b3;

        #200;
        key = 128'h009e_cb64_7744_f96e_37c7_935b_04d6_342d;
        state = 128'h14fa_9555_6aba_7fd4_9918_4cc6_9f2e_534a;

        #200;
        key = 128'h7d0c_b575_02f9_fff1_a70d_2e91_ff5f_1402;
        state = 128'h5408_ba07_6a57_c7c9_2ec2_7230_1d1e_e20f;

        #200;
        key = 128'h97bd_37f8_aadf_4293_a8e7_d7f6_c048_d04e;
        state = 128'h06de_76c1_320e_db4d_4c6c_e0f3_e36e_ddbd;

        #200;
        key = 128'h0c02_d387_dc93_626e_a3ce_514f_873b_054b;
        state = 128'h9956_aacc_bb42_4dbf_be18_82b8_2a6c_d395;

        #200;
        key = 128'h3fa5_3a69_40dd_0e6f_5bb9_e5e0_9e67_fa00;
        state = 128'h9bd5_9926_38a3_864e_83d7_fa2c_0813_dce2;

        #200;
        key = 128'h41d3_214d_3450_b33b_7f5a_5c74_d652_b732;
        state = 128'h4826_4ba5_f39f_cdd7_6d6c_cf6e_c858_8ba4;

        #200;
        key = 128'h706c_ceec_8031_b5bf_93b3_8125_7c66_7c1c;
        state = 128'hc930_f4a8_22da_1157_8b1d_bf3b_1d53_baa7;

        #200;
        key = 128'h6f22_427b_c56a_323e_26c4_eb95_f3a2_d076;
        state = 128'h013a_d705_c068_d592_be2a_7754_4e1a_dd35;

        #200;
        key = 128'h37c0_189c_942f_2385_206a_4c0d_a6d2_13f3;
        state = 128'ha691_e61c_5e2e_2338_a72c_0a12_cff3_be2a;

        #200;
        key = 128'he8aa_46d9_794f_472f_42c3_057d_a45d_560a;
        state = 128'h309b_ab2b_57ea_d356_e830_ce5c_1362_0d33;

        #200;
        key = 128'ha36d_3878_7748_e28e_d131_4613_a74b_83dd;
        state = 128'hc48e_2da3_c492_47d1_992e_dfbf_5f4e_7856;

        #200;
        key = 128'h1195_c949_883a_1494_22c5_8cff_1168_9927;
        state = 128'ha16e_8bf1_8c2a_b030_0ac4_d5de_df6a_91fa;

        #200;
        key = 128'h3764_ce93_7ddb_de8b_42c4_791e_ca52_5e96;
        state = 128'hd579_9f01_90ae_e14e_d441_585d_c854_072b;

        #200;
        key = 128'he172_8267_0fc4_793c_1475_e177_550b_fc21;
        state = 128'h24b5_407e_0b40_1260_0cdf_9061_1ff9_5180;

        #200;
        key = 128'haa0d_068b_2469_88d0_63b8_cc4a_aca6_8944;
        state = 128'h7e02_5130_b30e_63e0_e659_1afa_3aec_0c6a;

        #200;
        key = 128'h8431_2256_6191_bb92_6708_242d_028a_5df6;
        state = 128'h66e4_2821_2c98_53f4_f467_2728_358d_b17f;

        #200;
        key = 128'hffc4_35ae_4de0_45d5_7cf4_92a9_33fa_ca7a;
        state = 128'hc27f_f6df_3b4c_e217_70af_4192_a944_b11f;

        #200;
        key = 128'he833_6baa_b5f2_d712_befc_759d_ad81_6c09;
        state = 128'hfccd_bff6_4681_c91e_a8cf_6d37_532b_0c66;

        #200;
        key = 128'hc446_41af_d22f_d7c2_38cd_6aa8_a554_b843;
        state = 128'h6873_543a_1e5d_ef7f_73de_e3cf_a5e6_ed5f;

        #200;
        key = 128'hb788_3a53_c87f_b502_792d_59e5_0d01_cda4;
        state = 128'h1f0c_ecfb_6358_f56d_dc3f_f90e_597f_eb17;

        #200;
        key = 128'ha3c2_f711_7522_b02f_297d_90d9_af9d_2c12;
        state = 128'h4e9b_c4d0_11d8_0d07_7d01_3ba3_f5ce_a827;

        #200;
        key = 128'h7877_6e33_d1f2_e2eb_0474_0756_ef54_8aa5;
        state = 128'he529_3859_59b4_1e46_c346_c742_d9f5_e5c2;

        #200;
        key = 128'ha104_39d7_c789_958c_33a6_bfc4_42d6_1b6f;
        state = 128'h1abd_3a9a_2121_874c_839b_49df_c276_3fca;

        #200;
        key = 128'hfd7f_ab0e_6257_d495_7f52_73e5_7e90_473c;
        state = 128'h4f85_fbe1_ff7a_9b37_6513_355e_3040_023f;

        #200;
        key = 128'h5f9a_ce8f_6629_0faa_e3f3_ec56_52e3_1c39;
        state = 128'hc294_2807_db75_965b_bc5f_f5b9_5180_2e27;

        #200;
        key = 128'h497f_a562_b4a7_ad70_6e0f_2d97_e475_5c90;
        state = 128'h8a8d_59a2_08aa_2098_4d78_d64e_c49d_ab4a;

        #200;
        key = 128'ha6ff_734c_0325_2ce5_fd37_5284_e85b_5575;
        state = 128'he4a4_dd08_29d1_2452_769e_fd94_0dbc_6b7b;

        #200;
        key = 128'h9464_85a8_9d5d_ea20_efd0_4436_d51f_f33f;
        state = 128'hf520_2f6b_ebdf_5375_4381_33d0_a478_1fec;

        #200;
        key = 128'h739f_05c9_cf92_5322_0646_c7b3_f05e_0ad5;
        state = 128'hb96f_8187_e5bd_72c0_9c32_b055_ba30_f953;

        #200;
        key = 128'h9c3b_c24d_eaea_b6e9_a31c_900f_3443_3832;
        state = 128'h22a6_cf28_4a04_de87_0708_be9e_8df5_5559;

        #200;
        key = 128'h068e_a3c0_a5fe_a155_791d_3b8a_28df_7a40;
        state = 128'h0960_81fb_e4f4_2523_5961_0979_afae_099e;

        #200;
        key = 128'h5cbd_0535_06f5_20bb_1bd4_fbe0_c484_07ae;
        state = 128'ha894_0116_e396_1a68_2f97_9ca8_aa97_7eef;

        #200;
        key = 128'h3943_a994_5814_7514_9702_bda7_9189_6893;
        state = 128'h0eaa_498a_7b55_3461_3013_b3c1_a81a_eb52;

        #200;
        key = 128'hbb35_3c94_adc6_c7bd_2ec5_872a_9bd3_6768;
        state = 128'h55b9_3b24_4912_f4c4_2244_f6f2_a1dd_bec4;

        #200;
        key = 128'h4fef_b701_f3e8_5e5b_083f_e69e_082e_3d4f;
        state = 128'hae72_0242_a204_d871_b979_7fed_67e1_f08a;

        #200;
        key = 128'hdfa9_8e26_439f_2642_0a08_8138_3c89_5b48;
        state = 128'h8d2c_78b1_615b_12b7_9e30_b3ea_9727_0783;

        #200;
        key = 128'h257f_ba1c_81bc_1174_6bd8_d408_b081_b575;
        state = 128'hf152_d06b_e0f6_5cf3_a2f7_3d54_2151_09dc;

        #200;
        key = 128'hcbbc_bdbc_86da_ebbd_209c_db03_514d_c6ba;
        state = 128'h8ac3_09d3_f2fc_156c_5f32_b8ec_d4ff_e6e5;

        #200;
        key = 128'h989a_baf4_0811_4be3_d13f_19ea_0899_7f9d;
        state = 128'hc7db_e837_5998_4971_2a2a_3526_1d39_1de8;

        #200;
        key = 128'h525c_3df4_eb5c_ff06_9652_cd79_fe68_e2b2;
        state = 128'hd474_7b93_66fa_1c5a_5dbd_74ac_ffd4_d302;

        #200;
        key = 128'haa78_7977_5b6d_b296_2df3_0742_9c3d_d805;
        state = 128'h2455_722c_eede_0f09_fc80_090f_1c11_2ea6;

        #200;
        key = 128'h0207_98ed_49ee_abe0_ca8d_c5fa_091b_a7c2;
        state = 128'ha13b_23ea_b725_8c7b_0bc3_a492_a013_393b;

        #200;
        key = 128'hbd76_de11_0488_6aa0_f6b8_427e_deed_5f58;
        state = 128'hd1d6_fc34_8fd1_a29e_0469_67f9_6902_faa3;

        #200;
        key = 128'h7b9a_14d5_1f9f_e040_add6_e25e_b459_b331;
        state = 128'h54f9_b692_12f7_1f37_6c7e_98e2_03b3_7af5;

        #200;
        key = 128'h365c_39ab_5a4e_ae5f_0c8d_0f9d_4e41_5318;
        state = 128'hf7f6_fb27_98bc_f202_11ad_cf9a_16e6_beef;

        #200;
        key = 128'hdaf0_ad86_7a7e_0128_6054_ae21_5ffe_7c8a;
        state = 128'h6359_dd1f_8b39_1b4c_fbc2_2ab0_20ad_1188;

        #200;
        key = 128'h0381_b859_66c0_67fa_7891_958f_3bdd_1826;
        state = 128'h379f_6999_70ff_e5d4_6d6f_2062_7b7f_4d9b;

        #200;
        key = 128'h6be5_d501_ac0b_6717_d42d_6053_4df3_bacc;
        state = 128'h7758_0777_6927_4d4b_c735_06b2_47e8_06c0;

        #200;
        key = 128'had99_441e_4223_2b5d_cbc0_bde1_399a_3f85;
        state = 128'h8398_9aea_fc84_5795_aa59_aceb_1e7e_ace1;

        #200;
        key = 128'hdf6f_52ee_c226_e241_c67d_c2d6_e8ed_b68b;
        state = 128'hf8d6_03c4_c33f_1a6b_58db_cafc_ce18_e8e3;

        #200;
        key = 128'hc081_192e_4aec_43b3_7710_cd33_126b_a9b8;
        state = 128'hb281_8ecc_358f_3a9b_085c_6020_2042_e615;

        #200;
        key = 128'h5070_2a80_6519_5073_ebd5_e7eb_c2fd_57da;
        state = 128'h4660_a09e_d568_24e1_d8a3_fbdd_1fda_c44b;

        #200;
        key = 128'h3cc6_eb9a_f487_e775_793a_ee21_873b_4f6e;
        state = 128'h2795_e871_0f31_65eb_8b5d_0be5_263d_512c;

        #200;
        key = 128'h2b60_5ebb_0083_8737_68d8_43cf_e534_e9c3;
        state = 128'h3122_54c6_b957_1b1a_e19d_ab08_ce91_df99;

        #200;
        key = 128'h0058_1aa3_55ce_e463_fe43_06f2_0037_e997;
        state = 128'h6dd8_1d10_f57d_7e10_00ea_4ad2_a427_124d;

        #200;
        key = 128'h3ac7_2d7f_3159_fe3d_ada4_7047_9648_9c10;
        state = 128'hd3d2_6b7b_56eb_d7a9_bd25_ced9_91ec_52ed;

        #200;
        key = 128'hd547_a22b_022e_92ee_a07a_0c62_dad6_ce38;
        state = 128'h67ed_b810_f2ab_73f3_8c91_6402_1c37_1bb5;

        #200;
        key = 128'h6663_f497_84d4_814c_ba14_0df6_b6bf_53cf;
        state = 128'hcb2b_24bb_820d_463d_f7e7_9748_bf61_89a9;

        #200;
        key = 128'h69f9_95a5_4686_4830_f86b_47b0_3a31_2b8e;
        state = 128'h1581_1a88_3f92_ef8c_edbe_0b2a_37dd_61fe;

        #200;
        key = 128'hd3d9_b111_628d_8ddb_e5e6_3b10_af70_6ccc;
        state = 128'hd283_b853_c13f_0e85_8d9b_322b_08db_58e9;

        #200;
        key = 128'h9d1c_767e_db50_0903_88cc_736c_b020_7bae;
        state = 128'h11b4_5c6d_0ed6_0932_700f_df8d_19bd_3833;

        #200;
        key = 128'h8e42_07f8_2a22_4ed4_b19e_8a7c_7c17_f5c0;
        state = 128'h78ac_1a2f_b6d9_ada3_84b2_37a7_5aba_6acc;

        #200;
        key = 128'h27bc_9252_df29_0d4e_e01b_adda_6a61_4bac;
        state = 128'hb018_8a39_0c61_fba6_59bd_88b2_6ea5_b96a;

        #200;
        key = 128'h350d_80fb_3e87_5719_82cf_e1c2_78b1_02e9;
        state = 128'h45da_7ff0_d7f3_ee0a_6bd5_1454_1104_33b0;

        #200;
        key = 128'h0758_883b_f941_cf08_1327_4517_a89e_8814;
        state = 128'h88e7_f192_a534_5659_f9c8_71c3_99a7_623a;

        #200;
        key = 128'h3aca_c267_ffc3_e7e0_732f_f52b_333c_842e;
        state = 128'h3472_039e_83a9_6c84_4b32_6cee_7b2a_b395;

        #200;
        key = 128'h45d6_60bd_bcfe_16b2_258c_7d8d_7049_eb1d;
        state = 128'h5378_3955_e1ef_1cf0_e36d_db10_8fec_5f94;

        #200;
        key = 128'h23a9_6a75_3abe_dc57_ae56_fdb1_2bce_1cfb;
        state = 128'h2420_495c_80a4_e182_dd8e_7ece_3fbc_d167;

        #200;
        key = 128'h6cfc_1692_9faa_e02f_1c1b_428e_ad06_fb5b;
        state = 128'h9143_2189_a642_04d3_669b_b1ce_4436_bb4c;

        #200;
        key = 128'h0b0f_3da7_c877_f316_4795_b1ce_e529_a8dc;
        state = 128'he38b_58d0_7555_7fe5_3d04_334d_cb15_f2dc;

        #200;
        key = 128'h9d17_8f87_6797_86d1_5908_731a_b0b4_e6d7;
        state = 128'h063e_d61f_5927_a5e9_df28_597d_0fde_5860;

        #200;
        key = 128'h3f1a_691b_7348_81e3_7783_5717_5033_7973;
        state = 128'h237c_ceb7_52f1_3c44_6949_b3bc_24d2_06f8;

        #200;
        key = 128'h8f40_5347_8366_b4b5_0abb_e2a9_d610_f2f6;
        state = 128'h692c_1f97_4ea7_05cb_1f6d_a8a1_784a_d9b2;

        #200;
        key = 128'h5912_27e7_73da_4415_8487_384e_07e2_3a74;
        state = 128'h1b87_aa97_00c3_5cbb_1fa0_29a1_48da_fa44;

        #200;
        key = 128'h85a2_8bd0_b340_3311_d763_e49e_11ce_cac7;
        state = 128'hb964_a592_9048_a7d1_c740_6831_32d7_941f;

        #200;
        key = 128'h1948_0603_bbde_f705_8b4b_ff98_815d_80e7;
        state = 128'h5fea_2b7a_48ab_cfe3_7bbb_a3e0_0301_8b63;

        #200;
        key = 128'hcb20_3a19_1f5d_1608_ddde_9c9d_0eae_d9ce;
        state = 128'hd376_f258_1c8d_5090_560a_7712_ea3a_9d09;

        #200;
        key = 128'hb2b5_7ffb_affe_f5e5_be29_2ea6_cb04_cfff;
        state = 128'hd5aa_1433_fae3_5c6e_0ca5_97bb_0939_831a;

        #200;
        key = 128'h162a_5549_1030_83b3_7cb8_b042_83ab_5632;
        state = 128'hd077_35c5_e3e8_67ea_aeab_616e_a0ad_e2b0;

        #200;
        key = 128'h9735_f92d_9247_e805_3177_2ac4_7b2b_590f;
        state = 128'he431_ac35_fc9b_5aee_20c0_ee3d_917e_3015;

        #200;
        key = 128'h9fe4_e394_d24a_61b9_b5c7_c820_f2f3_c968;
        state = 128'h3b80_a4c0_e2d2_30b5_4362_216f_b832_fa78;

        #200;
        key = 128'hf808_655a_24e0_7f21_f593_05e7_ec83_0c4c;
        state = 128'hddec_5b84_f9f2_9f04_565c_7fc9_2126_9bf1;

        #200;
        key = 128'he840_8d1e_cd1e_8dcb_6e02_b800_51a3_c76b;
        state = 128'hbdb7_5727_631c_4fe0_f571_25ee_18b3_f7e3;

        #200;
        key = 128'hd389_4e48_ea18_a9c6_3bef_66c9_ec5f_d385;
        state = 128'hf0c9_b739_54b8_8415_2c2b_987b_acef_87cb;

        #200;
        key = 128'h1239_f9b4_1b4b_8131_6d93_4b4f_547c_8226;
        state = 128'he00c_fbb9_c499_2ce4_a04d_c4da_731c_7eb8;

        #200;
        key = 128'hb449_cfb2_cf85_6469_7149_d3bc_ff34_3ba2;
        state = 128'h00fa_df49_9f60_00bb_2e8c_e42a_7e46_90e8;

        #200;
        key = 128'h9a67_6c9f_b099_99fd_ef6a_6ad2_ee93_ad70;
        state = 128'h83fe_6bfc_a222_910b_788b_be73_1145_de4f;

        #200;
        key = 128'h1236_287f_6f78_aac0_8ae4_4aea_acf4_5424;
        state = 128'hda68_9f85_cfec_3c3c_0d88_607b_bcde_e8d6;

        #200;
        key = 128'hef7d_4a5f_1c40_50cf_51fc_90ff_fbb9_c841;
        state = 128'h2ecd_704c_de4d_dd4e_0c02_3be4_3943_79d7;

        #200;
        key = 128'h0d97_2f6a_dc76_ac3c_0428_48e3_7c8c_70e1;
        state = 128'h22cb_0f17_c1f3_852b_a97b_2c45_75d3_f726;

        #200;
        key = 128'h945b_8596_e666_edbe_6f92_adb3_57ed_7c1b;
        state = 128'h7def_d9b2_1725_17fd_adf7_3370_4981_0209;

        #200;
        key = 128'he906_e7e2_533d_1fea_8f87_3172_863f_e2e5;
        state = 128'h192a_c459_0899_c5ad_974f_92d7_4917_2215;

        #200;
        key = 128'h232d_7f79_81cd_59a2_b051_b475_9778_200e;
        state = 128'hb1a2_445d_e953_6b51_b35a_1f32_fe44_e0ef;

        #200;
        key = 128'haaa4_b223_c4e8_cf4c_0a01_c010_a99e_0d7f;
        state = 128'h85ef_695f_8cb3_ef19_4718_6b50_26dc_5e28;

        #200;
        key = 128'hf45c_b70b_c8c9_2af5_f10f_68b3_52ab_6c33;
        state = 128'h58ed_7e25_8092_6b9b_2f81_a1d2_2eb3_9a06;

        #200;
        key = 128'hf78e_b1f0_8be4_f848_c689_30c4_ab67_47e5;
        state = 128'h831d_8c76_9512_2106_2927_8ddc_03cd_05b0;

        #200;
        key = 128'h49d6_f0e5_5dab_ce64_93d8_cc91_ad28_41b4;
        state = 128'hc02c_50f3_4acd_4140_01e3_c7e1_5760_e6a1;

        #200;
        key = 128'h367c_a845_6867_7e4b_3b33_df62_2757_e279;
        state = 128'h6b4e_c724_2e8f_a8f7_68e0_2062_b068_9ead;

        #200;
        key = 128'h39c1_cc10_1659_d768_9e45_2ba8_3dd6_7c7f;
        state = 128'ha2f8_867c_115f_162c_0081_fa24_199c_f668;

        #200;
        key = 128'hbabf_94db_0fe1_5861_643f_534a_1f93_462b;
        state = 128'h2a85_886a_b528_3c5b_6222_79e7_2f99_2dcd;

        #200;
        key = 128'h05da_6dce_df8f_1e53_7c7f_cb4a_f631_8479;
        state = 128'hea9e_e356_2498_73f6_3982_bc3e_cc59_3794;

        #200;
        key = 128'h8918_ed5d_7c67_2716_fe90_0aa2_154d_cf45;
        state = 128'hb020_8a6f_9d1d_7438_65db_eba9_df28_885d;

        #200;
        key = 128'h2bfb_6ea5_5d57_4b5e_45ec_692f_60e2_e3e5;
        state = 128'h8b56_dbd1_395b_b197_b9da_f13b_46ef_defc;

        #200;
        key = 128'h3a91_3c09_5977_db98_b651_d984_61dc_52d2;
        state = 128'h8897_8acd_4ef6_c5c4_47c6_a36c_73de_c7f8;

        #200;
        key = 128'h8969_fd58_e77b_50c6_fbae_812f_a115_c064;
        state = 128'hd70c_c7bb_d28d_11f6_8d5f_62bc_5100_40b0;

        #200;
        key = 128'h53d7_d424_2ffa_9208_3fb4_a1fa_6468_dd29;
        state = 128'h9d13_d2e0_8c65_837d_0f11_9650_ea34_4b9e;

        #200;
        key = 128'hba05_ee64_125c_4f18_2eea_09e5_cd55_db24;
        state = 128'h101d_a352_99ab_711c_20eb_534a_af24_2ad9;

        #200;
        key = 128'h0160_e71d_cd8c_b51a_3d86_cf4d_a062_f36f;
        state = 128'hd6c3_325c_6b6d_5eff_3c9c_dc3b_bd1c_d14a;

        #200;
        key = 128'h8cd6_903b_db75_bdc1_2bb4_f616_f8e2_732d;
        state = 128'h9001_c39a_586d_2f0d_e071_3b12_dc5b_fc2b;

        #200;
        key = 128'hcae4_c700_34df_db2e_63fe_aeb5_3eb2_6a70;
        state = 128'h5818_e46b_efba_f4cc_34f3_da41_d329_e020;

        #200;
        key = 128'h0686_cfeb_838a_31b6_6df0_6e5a_8866_3ef3;
        state = 128'hcaa8_12df_e5c6_cd1e_f735_a7d1_4709_8b3f;

        #200;
        key = 128'h32da_8d39_e19b_3832_d0bc_91df_2470_decd;
        state = 128'h2dbf_e02d_cf0d_728c_4642_4974_8570_7bd1;

        #200;
        key = 128'h2219_d1a2_3698_1db9_cbd6_a996_5e90_a70e;
        state = 128'hd06a_2811_68c0_3ed2_f73e_e5d6_9eff_51f4;

        #200;
        key = 128'h3b8c_9f63_32df_ce1d_7485_a1e2_471e_ce18;
        state = 128'h5e42_8d4b_c76b_fc1e_4e6d_9f2c_4b17_5934;

        #200;
        key = 128'hb20f_02a5_47a6_38ad_2e79_97fd_0172_0c06;
        state = 128'hb677_2ef0_0631_e3d3_8137_90c3_3b8b_d364;

        #200;
        key = 128'h6835_a893_e1ac_b27d_bb7d_8b66_083e_10c5;
        state = 128'h2d01_a039_f4d5_898c_6bc7_da23_b87a_03b7;

        #200;
        key = 128'hac54_48d7_c125_37ff_a5fb_2f29_4de2_f1a0;
        state = 128'h0718_dfd5_a515_c9b3_4161_ce2a_c65a_2306;

        #200;
        key = 128'h735a_878e_c319_b9de_4b38_c592_4b4d_4767;
        state = 128'h3f75_55d6_30d4_42f8_96d2_5ad8_0750_2e4b;

        #200;
        key = 128'h8a54_7258_e684_b430_f74e_1bfa_627b_47fd;
        state = 128'h6e3b_1427_51c1_a1ea_9e12_2939_e0e8_c250;

        #200;
        key = 128'hd5d6_8979_8894_53c9_c807_ecdd_7458_db36;
        state = 128'h206c_f964_da92_546e_06e5_f419_df59_e1df;

        #200;
        key = 128'h66f4_0a4d_c071_804c_5574_7fff_7425_2074;
        state = 128'h7970_2ad3_7ee3_c9b8_31d7_42d5_c2d2_bdd6;

        #200;
        key = 128'hd9f3_693c_85b8_87a3_316b_6499_2bd7_d376;
        state = 128'hf35d_4f20_3f74_3deb_d27d_da40_cb90_59ca;

        #200;
        key = 128'h15b1_923e_1398_da24_7484_6d26_1d25_93e1;
        state = 128'h228e_aa3f_eefb_51cf_2e93_f4fd_5e77_838c;

        #200;
        key = 128'h361d_38b8_ef2b_44d7_e12b_12fe_23b7_c0dd;
        state = 128'hd43d_3dac_6d56_1e55_965c_89a6_d251_cb02;

        #200;
        key = 128'he4c8_5b40_7248_f275_ebcd_1cbe_188b_08e9;
        state = 128'h07b2_599b_6036_3024_32a4_0040_dbd4_8262;

        #200;
        key = 128'hc5d1_78df_bc7b_7efc_b0eb_daee_b306_2d50;
        state = 128'h8030_de88_89cc_448e_f18f_d556_ef79_7120;

        #200;
        key = 128'hc667_9be7_c24f_0382_ef72_2ef6_3fb4_5c0c;
        state = 128'h4f44_b2c7_22bb_3046_9adc_9870_64ae_ecfd;

        #200;
        key = 128'ha300_34db_3eab_7dbf_289b_af3e_346e_bcbc;
        state = 128'h3bbc_d197_2f18_3b30_8094_61d1_5e25_5817;

        #200;
        key = 128'h3a8d_b5ee_face_7113_34e5_7661_5caa_ea1a;
        state = 128'h3d96_b442_fdc8_5ce2_3f38_75e5_25a5_5969;

        #200;
        key = 128'h9472_6f78_b923_8598_a171_f2ac_d289_c6d6;
        state = 128'h17f8_d14e_c665_3034_8c06_ee08_41fc_e005;

        #200;
        key = 128'h9d88_54c7_7765_d7c1_564f_ab7a_c207_d8e5;
        state = 128'hfb2f_4d2c_476d_212e_20ce_a5f7_2b28_25e0;

        #200;
        key = 128'he2fe_4840_8236_2712_6a6d_18d2_fda2_6c95;
        state = 128'hce9f_5559_8c74_8558_1acd_ab88_31ae_37eb;

        #200;
        key = 128'hc634_374b_7fb5_f707_942f_e648_2a2b_4006;
        state = 128'ha5ef_8a13_773e_97f6_7be8_ead1_6c8b_83c4;

        #200;
        key = 128'h816d_091d_c65e_3d67_75bd_4493_c8b2_3e3b;
        state = 128'h2843_915f_84f4_1fc1_c59e_6edb_da9a_969f;

        #200;
        key = 128'hfb50_f396_1bce_5ab8_3b89_f67c_7a38_0cdb;
        state = 128'h4285_04c1_c8ff_b5db_4674_c22a_a2c3_1b06;

        #200;
        key = 128'h1cfc_a925_8f8e_1ecd_9fe9_39ae_5004_4faf;
        state = 128'h0535_0cf9_a159_d030_6c37_77c8_a41f_92cd;

        #200;
        key = 128'h69f5_0037_c0a6_64f3_d854_3392_bfcc_b81e;
        state = 128'hf566_3e88_5d6c_623f_4c88_e41f_ac7a_1797;

        #200;
        key = 128'h2532_2cf2_5744_9bfb_7ff9_ccae_01d2_c848;
        state = 128'h075a_a732_ae6e_4600_65e9_9464_9cd6_c7c5;

        #200;
        key = 128'h04ba_d8b7_479e_0b7b_c7d7_a8ed_1ba5_5dde;
        state = 128'hef50_92f2_7605_dab9_a7ef_3ed8_13d4_29d6;

        #200;
        key = 128'h5631_6723_ec16_887f_1714_4772_d052_1090;
        state = 128'hc662_184d_ee1c_fe10_6f15_7430_bebb_1719;

        #200;
        key = 128'h6e69_65cc_b2bc_10d3_f976_8637_65a7_d6c0;
        state = 128'h05cb_4e78_a322_6cf2_35f9_357e_689b_b381;

        #200;
        key = 128'h6553_2c5e_0da5_8384_0677_6ab9_82d7_6005;
        state = 128'h3bd5_2187_2535_3a8f_4980_ee04_a578_3317;

        #200;
        key = 128'h37ee_0cff_e2c9_42d8_dd19_867e_4400_4b10;
        state = 128'hd587_78c0_1560_a1f0_40c1_3a64_0f2c_a9d7;

        #200;
        key = 128'h86a0_d241_8e04_3cc7_de7e_07a8_be24_870f;
        state = 128'hb6d2_aca3_9b6d_5ad8_ea58_0f44_11ea_9a4e;

        #200;
        key = 128'h589c_89c3_e624_7f69_25e6_f96d_f53b_f60b;
        state = 128'haf9a_f5e8_9c02_7e4b_6cf5_8633_b591_4bc6;

        #200;
        key = 128'h4145_245f_8af2_9091_0894_1a63_1521_fb36;
        state = 128'h98a3_5370_8aa2_0348_4b7a_7e09_2974_3442;

        #200;
        key = 128'hd490_9ba0_c434_c9e0_147f_9acb_f696_ee3c;
        state = 128'h8429_8cf6_f3d3_2a08_4a1c_b671_7d29_f0be;

        #200;
        key = 128'hd0c7_74ca_ccc4_fd69_4d87_be5a_766d_5e98;
        state = 128'h8834_e5c1_4dce_c500_31ec_3caf_e0d7_62aa;

        #200;
        key = 128'hd51a_992c_dafb_b99e_21c6_bfc9_8f7f_b736;
        state = 128'h0f82_fc82_c4f3_3dd4_3158_fbd2_9361_a2fe;

        #200;
        key = 128'h6629_0de7_3c5a_3fbe_a7ec_a226_ca7f_f9a4;
        state = 128'h0bd4_2729_bfdf_2668_322c_61bb_e1a8_5072;

        #200;
        key = 128'h57d3_8d25_bbd2_dfa3_e1c1_5def_173a_1274;
        state = 128'h0c75_01b7_4912_b721_6351_4df2_4850_fa60;

        #200;
        key = 128'h97a2_565e_e4cc_87ce_ef65_89d9_6026_6f6f;
        state = 128'h56ba_c568_2fbe_0cd8_2378_00da_0a2f_de1d;

        #200;
        key = 128'h406b_4bde_cd75_a8c4_1b9e_ecb1_35a6_9b1b;
        state = 128'hb2ea_6ade_75f8_390b_3c97_4b6a_712f_f62b;

        #200;
        key = 128'h4323_5eee_ed3c_3d59_a4f8_7a70_977c_d8bb;
        state = 128'h8c5c_b926_0a7b_eb02_f8ad_1176_0f3b_2091;

        #200;
        key = 128'h6060_1602_5d5a_ff11_8ebc_bc25_ceda_866d;
        state = 128'h1aae_a5bb_dbb2_f8ef_d094_c010_bd4b_387a;

        #200;
        key = 128'h8336_e0b6_3115_e56d_e282_1ff9_0416_ec67;
        state = 128'h64d9_b500_e918_b73e_ab65_98e5_6025_e828;

        #200;
        key = 128'h203f_92a7_40a0_7853_97fb_078f_5444_41d1;
        state = 128'hee17_45c4_66ee_6301_2d1f_0766_6bdd_eb26;

        #200;
        key = 128'h5136_a93d_40ee_5b17_387c_d679_6486_f48a;
        state = 128'h190a_1cfc_68df_88b9_9fea_6b73_708f_8573;

        #200;
        key = 128'h5578_c93e_4c00_f6d3_5d57_72d4_3573_82b9;
        state = 128'ha574_7c78_fc14_1000_e503_778a_253d_9205;

        #200;
        key = 128'h5285_f75b_d1b0_1da4_3e98_929f_22ed_3a96;
        state = 128'h87cf_5dc1_cd38_193f_8004_8a34_47ff_4862;

        #200;
        key = 128'h7c76_331e_4eb1_e1c0_4c7b_aff2_9c20_6105;
        state = 128'h5cc1_815c_d6bb_2e83_35ac_49cd_5ef7_2ac6;

        #200;
        key = 128'h9df5_6907_a7f3_3821_b7b7_2024_3995_764a;
        state = 128'h8f38_0e83_a66d_6293_866f_e79e_c4ba_f251;

        #200;
        key = 128'hee72_b98d_b8b6_f0ee_9cf5_b288_08e1_a52f;
        state = 128'h7b04_3763_8bb5_5eb1_6175_923c_eaec_5d6e;

        #200;
        key = 128'hc5bc_9ae4_5f0c_683b_68f7_7691_763a_7071;
        state = 128'haf65_6e6e_7ca8_9b91_172c_d262_6f44_aba6;

        #200;
        key = 128'h12ba_09dc_6e4e_fdf0_bb18_20eb_7674_64ff;
        state = 128'h0323_22fd_0b90_de9b_7846_14ea_b10d_6645;

        #200;
        key = 128'ha44c_f44a_4913_a845_3a7e_edbf_27d3_5515;
        state = 128'h0acd_e707_0de3_9360_7b6e_6c98_f462_b3af;

        #200;
        key = 128'hb2a1_4b81_5049_7ffa_619a_42e3_f517_c8d1;
        state = 128'h228b_7f22_527b_7d7d_695c_8d3f_d845_f045;

        #200;
        key = 128'h2a6b_b7f7_a4c5_9676_265b_6713_e1e5_69eb;
        state = 128'hb820_1f31_fb45_dfa5_a06b_7ff0_d611_5456;

        #200;
        key = 128'h0619_99cf_183a_8459_aa07_ecf7_255e_6691;
        state = 128'hc5a7_0e8e_4116_118b_a375_2d20_8df0_0613;

        #200;
        key = 128'h809b_e781_8331_8009_53ee_63fc_7463_27d4;
        state = 128'h1a70_2af6_296e_eb25_e61d_fd49_519e_15b3;

        #200;
        key = 128'h60d4_a739_42fe_01a3_bbd4_e282_b3bc_4901;
        state = 128'h9a27_177d_06dd_8eb1_24cc_4701_0c6f_a227;

        #200;
        key = 128'hb5ed_7f8c_9336_c9f3_17e9_fe3b_99be_55e2;
        state = 128'h03ae_70b4_53a5_02fe_f24f_bd1a_f41f_0422;

        #200;
        key = 128'h1c6a_cc40_028f_4fe0_4d1e_9efe_3311_2272;
        state = 128'hcd1c_b2d8_4d26_c933_aa84_c37a_d4b1_1915;

        #200;
        key = 128'h9de3_f694_c960_83fb_0ec0_67d1_f13a_9d7d;
        state = 128'h7c47_0d83_7c0b_425b_9d11_cc54_e0ff_17a7;

        #200;
        key = 128'he2f5_e985_7041_aee8_c624_0506_b6bf_c46e;
        state = 128'h6304_b032_0d27_2fef_f982_849a_4e9d_48f2;

        #200;
        key = 128'ha026_bb1a_e241_e7b8_5f01_45c1_5379_d896;
        state = 128'h84df_d5c0_b423_7a2e_2fe8_cef1_a969_488b;

        #200;
        key = 128'h1cf7_0858_1348_21c5_4a42_0fc4_807b_34d1;
        state = 128'h3286_a500_e250_7eb6_1eba_05c4_7de2_0a71;

        #200;
        key = 128'h8509_5e3d_b042_485b_e977_90ef_4d58_c8a4;
        state = 128'he857_f1eb_1566_fac0_3b88_c76b_cfbb_d532;

        #200;
        key = 128'h148f_f82d_b70b_9460_d0cc_133b_6733_820b;
        state = 128'h520b_fe40_97ea_bcca_25a1_6914_267d_0134;

        #200;
        key = 128'hf398_db4b_c66b_f26a_62b2_3d98_c5c4_3453;
        state = 128'hdfcc_9dbc_d146_a534_2d10_1a51_2e8f_9c3a;

        #200;
        key = 128'hff7a_a2cd_dbcb_53a5_58a7_c1f7_a950_707d;
        state = 128'h813d_491b_f9b6_a84c_4759_5e05_4ebf_1661;

        #200;
        key = 128'h333f_c411_aa41_56a1_2667_e278_1d3c_391b;
        state = 128'h6950_1acf_35bf_6759_1db0_52c8_d8d5_e471;

        #200;
        key = 128'h3870_2d3e_9ae1_568f_3d57_a3e7_a03e_8b21;
        state = 128'haf17_6009_214b_0139_7fef_b82a_1ddd_af22;

        #200;
        key = 128'hd344_51c6_29c7_9365_8215_9d17_31d6_7fd3;
        state = 128'h2368_4e88_6e71_d88d_6e7c_c80a_1f12_fb98;

        #200;
        key = 128'h7bec_cfcf_db99_9032_9a14_b109_6212_8139;
        state = 128'hd151_8151_2409_6eba_eba0_66bf_5a88_deff;

        #200;
        key = 128'h4311_839e_9780_24f0_e9d6_5aa6_687f_2c63;
        state = 128'h7404_4a2f_8137_b7ba_7482_16d6_d911_32be;

        #200;
        key = 128'hc5d9_10c8_db95_2cc5_c066_6905_ba52_30e8;
        state = 128'hb378_8e5e_daac_9c5f_2d65_ff00_e41d_a037;

        #200;
        key = 128'hc547_3eb4_5704_ebc1_8d6d_897e_eac9_913f;
        state = 128'hdc24_ec88_2579_add0_cc90_3d5b_ee8c_cc88;

        #200;
        key = 128'h842e_4fe9_c9c7_279e_d122_93ce_98a5_11cc;
        state = 128'h5bb4_b39c_bb43_9ed7_74fd_ea9f_4c23_18b2;

        #200;
        key = 128'hbb58_7872_8379_e910_f5f3_2bed_bdab_ba9d;
        state = 128'hffc8_fbd5_fa42_b2fd_aabb_765c_e3c6_106d;

        #200;
        key = 128'h0105_c9cf_e847_bfd0_5430_6df5_b2e8_b33c;
        state = 128'h2460_6911_4fda_ed3a_37c6_e925_d1d3_548c;

        #200;
        key = 128'hb68d_7ee4_fb1d_1073_3b0e_19a1_f34b_bd6d;
        state = 128'hb465_7cd3_5272_6263_7ae5_ea09_bc38_87fc;

        #200;
        key = 128'hc29a_e0cb_8276_471c_c883_2e1b_8e6d_3eba;
        state = 128'h34c4_d7f0_5e09_2746_b5de_3a28_f17b_4e49;

        #200;
        key = 128'h69e0_5723_759c_da93_86b4_0610_5719_d003;
        state = 128'ha4a6_3dbc_1a2b_a81a_6b72_ec24_33c9_f6d3;

        #200;
        key = 128'h3376_6445_8456_ee7e_757d_3e8d_f683_ea4a;
        state = 128'hab32_45c0_bbbc_6f08_f2a7_c12c_9a0f_8baf;

        #200;
        key = 128'h0835_df51_8ddc_2edb_9aa2_e0fd_bd49_2fcd;
        state = 128'hb925_b1ed_ff5c_fcd0_7a02_9b83_9034_b532;

        #200;
        key = 128'h1ada_33b6_38ec_7ac0_9746_742e_005a_7af5;
        state = 128'h7c7e_9227_09fc_f9d0_c466_1eec_dd0a_928a;

        #200;
        key = 128'he303_e5d4_2abc_7b4a_e262_f61f_5e57_7993;
        state = 128'h2c08_a245_f360_6427_f02c_3ce4_49cf_9dee;

        #200;
        key = 128'h7581_499e_0c70_66d1_41f8_8d84_1ac1_06d6;
        state = 128'h1868_067a_3077_7eab_7911_cf7d_e722_a20c;

        #200;
        key = 128'h3222_3a0f_5767_95bc_1409_2dcc_602c_2bce;
        state = 128'h1d9c_1c7e_6a64_4c2e_51ba_c52a_ec79_ab91;

        #200;
        key = 128'h8593_0ff6_ebff_5ded_3ccd_1f9e_aa11_8ab8;
        state = 128'h0f28_b6fd_ec2d_c9a1_031c_5a13_68dc_6285;

        #200;
        key = 128'hbafa_2edb_bffa_5a21_b928_70b1_9612_93c2;
        state = 128'h1af8_8013_78c2_fd7c_8346_f83c_e5da_477c;

        #200;
        key = 128'hb1e4_6f3a_78c7_dbca_7654_10b4_5c77_6631;
        state = 128'h206a_66fe_7347_ec43_a725_3ef1_cde5_653b;

        #200;
        key = 128'h3c0f_2b3a_365d_0fa6_67e3_8b94_2e23_feb2;
        state = 128'h7767_c957_1c2c_591e_e68f_7604_71b4_b561;

        #200;
        key = 128'h5f5a_ea99_e397_a3b7_df22_fb53_edb3_2ec4;
        state = 128'h167e_f143_09b2_c1b5_9663_7dbe_275f_e297;

        #200;
        key = 128'h8b4d_3694_ebdc_d07c_4e28_eadf_c839_9fdd;
        state = 128'h0f79_dfec_4705_ff9e_b1e9_07fa_22a7_5163;

        #200;
        key = 128'hb658_687d_2b25_8b85_7ea0_4ce6_c189_dfc5;
        state = 128'haef1_94b4_9a89_04a1_1496_251e_1799_5e40;

        #200;
        key = 128'h4a21_db1e_fe92_6c06_c128_2255_f799_3de3;
        state = 128'hb85c_82fd_5dd5_4461_9dfe_5262_9712_ec7b;

        #200;
        key = 128'hcad8_5515_5103_eba1_b02c_fa09_a138_0631;
        state = 128'hda37_20ac_82c7_fcee_7067_6dfe_6407_aaa4;

        #200;
        key = 128'h9ebd_e7f8_3a24_0472_5953_8454_bd57_2325;
        state = 128'h31cf_357f_76b6_46f3_d5ac_5d32_7e51_ded5;

        #200;
        key = 128'h6e8b_7906_550b_63b5_a151_ce46_8c3f_76cd;
        state = 128'h1c0a_1a32_5e8e_8dfd_af31_ac9c_c960_5683;

        #200;
        key = 128'hba5a_b614_8cb6_9299_b395_5578_fea8_d308;
        state = 128'h83ee_5f14_18c0_7751_38eb_087e_bd72_3f48;

        #200;
        key = 128'hbd3b_aec0_c775_468a_1ca4_4eed_d821_8927;
        state = 128'he76c_33b0_a0bd_779f_b63d_26e1_5c68_9883;

        #200;
        key = 128'hd724_04a5_9c63_fbef_9530_ba39_4426_7988;
        state = 128'hb2ac_eafc_c8bd_f7d6_54b1_489f_4701_79df;

        #200;
        key = 128'ha80d_3a92_98a5_4ca1_6e72_7de8_420d_eefd;
        state = 128'ha214_b610_528d_a47d_49dd_0af4_3243_a067;

        #200;
        key = 128'h0f98_5cb2_a135_d219_2712_ce34_1a6f_acdf;
        state = 128'he53d_bf87_935b_1ddb_5a2a_9a2f_04fc_0196;

        #200;
        key = 128'h534e_1010_5656_d248_0dc7_2aec_bc67_fa82;
        state = 128'h5cff_335e_162c_a645_1245_3fb9_0214_70af;

        #200;
        key = 128'h0800_8de7_f09b_ba3b_5326_36a3_c833_9436;
        state = 128'h20c0_a229_72e4_9494_9794_da2d_7360_96e0;

        #200;
        key = 128'h668f_7935_718f_f482_f07c_6dc3_5f70_c65d;
        state = 128'hfb0b_eed0_eb3a_0572_5a7c_3dd9_612d_7e6a;

        #200;
        key = 128'hfe2b_9e15_1246_ee74_20f8_d81a_d073_12dd;
        state = 128'h7865_d6af_3092_b11e_d216_a1c3_02e4_d3c5;

        #200;
        key = 128'he952_b5a6_71b6_3044_b381_97a6_7474_848a;
        state = 128'h98b3_5e91_127c_e929_29fd_66a6_a3e1_015c;

        #200;
        key = 128'hd6cf_7a2d_343d_569c_fe7c_bbbc_d6a6_5c56;
        state = 128'hdd7a_c5b5_0368_9f53_64cb_8281_e0a0_0513;

        #200;
        key = 128'h6193_d2fc_a332_96d4_bb15_5302_8a80_35f4;
        state = 128'h9397_4c9e_1b31_41aa_ce93_0e2d_4ef8_0ffb;

        #200;
        key = 128'h15a3_93b1_6ea7_31e8_ef30_ee60_d531_c82d;
        state = 128'hbef4_9a9c_a9d3_a82a_e640_4e57_93d2_d71d;

        #200;
        key = 128'h1b9a_1988_0fd3_d41d_161c_101c_b7d3_fc01;
        state = 128'h0201_5a0f_a568_62d1_600f_951e_0ec1_8d3b;

        #200;
        key = 128'h08fa_2cef_5802_0c69_7bbf_864c_5455_4940;
        state = 128'hcecd_61ee_bc1a_7e4f_65e4_b75b_089a_5141;

        #200;
        key = 128'hb69c_a195_25d8_b40b_e678_9fc9_57da_b3d5;
        state = 128'h3852_6abb_6825_ba12_41e4_e130_492e_8623;

        #200;
        key = 128'h8a16_4424_c3d5_708f_6601_5878_4e4e_ec24;
        state = 128'hd59b_0643_3ea5_c6b1_32a2_46fb_c835_e89c;

        #200;
        key = 128'hb0dc_1ec6_cfe4_cb73_4770_0808_598b_1816;
        state = 128'h361d_8ff8_2579_de9e_735b_af4c_ae2d_c1dc;

        #200;
        key = 128'ha1d4_6d63_4764_3a72_0af0_b494_4841_7e97;
        state = 128'hf8d3_0854_765e_7eef_a543_74cd_e024_b5bf;

        #200;
        key = 128'h6a48_9ee7_6853_1de0_6660_17be_d3ab_8772;
        state = 128'hb78b_cf88_1f51_e0e8_9789_1bbd_8a9f_c7f3;

        #200;
        key = 128'h399d_8a10_2407_1483_1591_7437_88ca_c9a1;
        state = 128'hadf8_568a_4432_8abc_e7bd_cc08_edbd_bbd5;

        #200;
        key = 128'h029b_0704_0571_d4fe_388d_90a4_adbc_195e;
        state = 128'h3515_2310_35a6_c650_f2aa_efb2_eca7_13a5;

        #200;
        key = 128'h3b92_a7d8_a663_8b96_2ef1_ce23_40c2_d646;
        state = 128'hb7ba_cadd_a7a4_a799_9587_e940_98e8_9492;

        #200;
        key = 128'h72ff_f710_f023_e59c_71e4_d3f9_e1c5_93af;
        state = 128'h7ec3_8e0f_4cc0_5b16_d98a_cca5_80c2_fd9f;

        #200;
        key = 128'hfe72_7371_21df_2524_105e_b88a_bee4_8f73;
        state = 128'h307f_7da7_d83c_4617_fd32_ef84_31aa_79ee;

        #200;
        key = 128'hd4b2_b499_c79f_81bf_87af_8da1_86d1_e0c9;
        state = 128'hbfb9_0c9a_dd47_ff47_46e1_9e9a_c001_ae54;

        #200;
        key = 128'hf226_63b1_802e_97b4_e5a5_16b9_896e_19d5;
        state = 128'h24b6_284f_bc86_7463_0ca3_f9c0_47a3_9356;

        #200;
        key = 128'h305e_c0e8_f70b_546a_e502_19af_3b57_9f0d;
        state = 128'hd6b4_1342_bc10_136a_51d9_b930_8d14_30ab;

        #200;
        key = 128'h8660_3427_09a3_e21a_f65e_b37b_d455_2131;
        state = 128'h8293_caae_de4d_ff48_ebb1_75df_c83f_26a6;

        #200;
        key = 128'h1778_9f94_09ae_ba1d_17cb_77b8_8d70_f8f6;
        state = 128'h2fba_5fea_0e76_0429_fed0_ad8e_111f_1107;

        #200;
        key = 128'hc9b5_6141_2dd5_b6b5_7528_a5dc_dcb0_9b47;
        state = 128'h4d94_e6f5_612f_3cdf_0283_c7a3_e84d_f04a;

        #200;
        key = 128'h25a5_3fe0_00b7_438c_f3e7_7fc8_b1bf_0140;
        state = 128'he35b_cbcb_2b6a_c9b2_347f_3720_0047_8fae;

        #200;
        key = 128'h45a2_1478_8889_bd95_9eb9_c4eb_dc9d_0839;
        state = 128'h714d_7187_d4f5_d889_c8c3_e3e6_fe33_587c;

        #200;
        key = 128'h4d85_7d30_dc52_801a_4bb3_a0ea_2daf_689f;
        state = 128'h40c7_a180_8365_1f07_0530_4a8a_c5f3_cc34;

        #200;
        key = 128'hf303_1003_dd7f_9593_da82_4f8d_24cc_7b4d;
        state = 128'he907_3fb5_d196_5873_e304_d066_320e_5bcb;

        #200;
        key = 128'h10e5_51e7_de48_c55a_f480_cfa7_eb4d_c7d4;
        state = 128'h3536_5aaf_a43b_2524_4cdd_b3d4_9324_ccd8;

        #200;
        key = 128'hd182_df80_f03a_03ae_6f81_b948_4338_a893;
        state = 128'hb4b4_d20a_5d7b_b6ef_204e_e86a_e904_fd28;

        #200;
        key = 128'h43d9_57f1_00df_1ce6_e32b_d163_42e8_046c;
        state = 128'h7ac6_6743_c017_78a5_30af_ba03_2b1b_b011;

        #200;
        key = 128'h90d8_6810_d9d9_a69e_8676_12b6_cdd9_ec84;
        state = 128'h598b_f5b6_3d60_21b6_968a_b4f6_90c1_dc1f;

        #200;
        key = 128'hc200_987f_b6d2_5850_9384_f8d8_1005_d9d4;
        state = 128'hecab_999a_0e13_aa8e_e3c5_a613_bc75_65a3;

        #200;
        key = 128'h003b_9abe_ffe5_d089_d3e9_f148_2aa0_89e6;
        state = 128'hfcad_3e46_a1f4_b2ab_afff_5fe0_431b_b95b;

        #200;
        key = 128'h9675_b39e_2a91_cd79_fd6e_ff66_3fbf_ee9a;
        state = 128'h3056_823d_c0fa_0686_c3de_ae73_d5ee_7913;

        #200;
        key = 128'he1ce_ca16_4eb8_ce22_0607_7285_ab32_708b;
        state = 128'ha8e6_f87e_ca5d_e6e1_eaef_48ed_6e6b_c0f0;

        #200;
        key = 128'h32c2_4859_5735_a1a3_8672_4b01_1b5e_a9e2;
        state = 128'hc06e_c461_2634_dbb1_d80c_12a6_ce46_1fc7;

        #200;
        key = 128'hd0b1_ef6e_9089_84cf_9185_f843_a494_843a;
        state = 128'heb2f_4efa_e708_348a_4700_fa46_05f8_7564;

        #200;
        key = 128'hbdb6_1ef3_3476_7d79_9efb_fdac_512d_ae49;
        state = 128'hb5ce_e18e_4863_988e_2664_6244_20cb_dda6;

        #200;
        key = 128'h5595_1f8e_f90c_d8d5_1c43_ae58_c450_2dd8;
        state = 128'h4231_1258_2fab_c806_1117_2811_f454_c63e;

        #200;
        key = 128'hf33f_7a35_fad2_c62b_eb9c_f646_6f9b_48b4;
        state = 128'h40a6_1b9c_7f79_bbb9_f99e_def5_b378_d4b9;

        #200;
        key = 128'ha9de_cbfd_181f_b2de_241b_89dd_57eb_b7aa;
        state = 128'h970c_92ef_727d_ef7c_205b_612b_6435_f9ee;

        #200;
        key = 128'h05cb_b901_518e_f91a_605c_2c4f_159d_4de9;
        state = 128'h4069_4c6a_478e_1c5f_f724_bb8b_d20c_514e;

        #200;
        key = 128'h3b19_59bc_dfd3_2131_04c8_a7ce_a152_ab9d;
        state = 128'h816e_6b4c_9b26_564d_a99d_6c9a_09f4_c9e6;

        #200;
        key = 128'h4eec_6a5f_992d_96b3_22af_d716_c497_c4e9;
        state = 128'h1d4d_fa2e_120d_f387_2bc1_e52c_2823_10a8;

        #200;
        key = 128'h8d49_4c6a_b868_b2d3_41b9_2f52_b85a_2d01;
        state = 128'h70a6_5ea4_9fc2_6d7f_3da2_c60a_7213_ef6f;

        #200;
        key = 128'h6917_7d59_5cb9_d5bb_75e3_72a7_ff53_194f;
        state = 128'h8a70_05dc_e372_b8c1_1289_be60_73fb_f4fc;

        #200;
        key = 128'he0c2_4c62_c59c_6d35_89e5_178d_ebef_0aa9;
        state = 128'haa1d_c318_2e15_677b_439b_0651_86cd_fadb;

        #200;
        key = 128'hfc87_7304_27d6_d7f8_6cb0_1717_a5d1_72c7;
        state = 128'h6525_fc17_52a5_2187_85e5_8481_b6aa_16c2;

        #200;
        key = 128'hb49b_2147_efa8_b25f_be4c_896a_0009_4f0c;
        state = 128'h6658_c079_5165_049f_d39d_1fec_1f22_7b5e;

        #200;
        key = 128'h795d_eec5_870f_bee0_6a83_1df0_e3c3_8cb1;
        state = 128'hbbc6_2a72_97d2_4b33_c147_81cb_585b_6e17;

        #200;
        key = 128'he461_d1ce_0490_58d2_c323_7951_5005_5569;
        state = 128'hdb24_d3f1_74bb_6029_edc4_1237_c1f0_279d;

        #200;
        key = 128'hc25a_62b6_5d36_a8f8_f4a4_ed62_4a66_e02f;
        state = 128'h7e52_6173_e2c4_4771_b236_b85f_bbde_1284;

        #200;
        key = 128'hc0ea_7aa6_619e_e483_52d0_2c10_2016_28ec;
        state = 128'h1aed_41db_7a99_2aed_57f7_b4ca_dcb6_f926;

        #200;
        key = 128'h41df_0a63_73aa_429a_9fde_eab8_1fd7_229a;
        state = 128'h608f_d7bd_3ed8_8fd7_3df2_442c_3dfa_a285;

        #200;
        key = 128'hb6ba_7ae0_d442_5ffa_1ed4_d8a2_8efd_bdcb;
        state = 128'h4b8c_5704_4b3d_70cf_5b5b_749b_51f7_5084;

        #200;
        key = 128'hdc14_94e0_78c1_88e8_9cb5_62da_6016_8a5b;
        state = 128'hb043_ee2a_fbdc_c177_07c9_8173_966f_b5a7;

        #200;
        key = 128'h4882_c748_40cd_8db7_9175_224b_7444_1d48;
        state = 128'hcd8d_092c_a6be_168b_379d_918d_6b52_ccc3;

        #200;
        key = 128'h226d_8711_d531_163a_c2e8_ad98_5132_f1f8;
        state = 128'h194f_e0ef_446a_7eee_e8bc_7aab_5774_44af;

        #200;
        key = 128'hf982_8538_9d66_04bb_810a_a87f_f803_e0aa;
        state = 128'hf180_b16e_d4d8_c07c_49ee_ce20_e0fb_6110;

        #200;
        key = 128'h761e_307d_1a62_601e_f59a_4378_b5a8_03de;
        state = 128'h512f_854e_583a_f9b7_6348_6991_b432_a496;

        #200;
        key = 128'h2e20_e692_516b_e11f_8f58_a03c_0ad2_9701;
        state = 128'h6b76_deba_725b_4f03_508a_2675_3bd0_ae8e;

        #200;
        key = 128'h5b66_d7c6_56cb_446a_c112_a49b_84ef_c8a7;
        state = 128'h937b_c28b_46af_e1be_053a_ba7a_1a27_1e4d;

        #200;
        key = 128'h1230_4600_bc9b_7259_de5d_9ce2_3ab4_89df;
        state = 128'h1956_7605_2de4_f25f_990d_5185_c22b_bb1c;

        #200;
        key = 128'hbe03_19bc_c1d9_8097_ef1e_1123_8d84_7e63;
        state = 128'h004b_7f2f_e2f2_f948_60dd_5c1d_5942_6399;

        #200;
        key = 128'h96e4_becc_71e2_4462_3e28_2298_db6e_0c5c;
        state = 128'hf3e2_3ce3_461e_a5b7_b2a7_5eb8_907f_3a3b;

        #200;
        key = 128'hb9ca_3d6b_2f96_2bd4_3119_c248_cd48_a99d;
        state = 128'hbf07_9500_7168_f179_3891_7dbb_1bf2_ab9e;

        #200;
        key = 128'hfdef_7d38_4cf4_0eda_b585_2c05_5606_3951;
        state = 128'hcb87_12c4_253c_ff69_14bc_e0f6_b055_8062;

        #200;
        key = 128'hbfba_4628_e23c_b28a_b6e4_bc06_daa4_11e3;
        state = 128'h18f2_7d4e_5b79_1e12_08a8_53ab_81e1_8473;

        #200;
        key = 128'hd246_b6c5_98be_5da9_a978_02a0_efdf_8e1b;
        state = 128'hc35f_bade_0010_cee2_f2be_21f2_4106_6d9f;

        #200;
        key = 128'h5388_eaf7_78b5_03d4_73a9_2614_a250_1a37;
        state = 128'h70ac_cbec_be6a_b0e6_f8e4_cbe4_40cc_7f24;

        #200;
        key = 128'hc87c_f705_699a_d7d3_1339_af76_5481_060b;
        state = 128'h8934_1787_d6f1_92a2_a343_1c48_f854_b3eb;

        #200;
        key = 128'hafad_0951_caff_1052_2800_6870_1dbf_b2df;
        state = 128'hc48a_b23c_d0e4_6094_42c7_f196_6543_e3c1;

        #200;
        key = 128'hb1c4_977a_1cb7_c65b_7eec_ee4b_641f_22dd;
        state = 128'hed97_f6a9_d335_4871_373f_2902_ebce_2d32;

        #200;
        key = 128'hd65e_f162_36dc_9148_404a_29d5_fbc2_e667;
        state = 128'h1273_ac5d_87dd_4ffa_26af_2542_fad4_a907;

        #200;
        key = 128'h47d5_d651_3b57_48c6_744b_4ca6_60ba_b8fa;
        state = 128'h1e06_725a_9cb2_eb0c_80cd_a463_90d3_f175;

        #200;
        key = 128'h5d2f_e463_6fc2_7820_1b27_9068_5775_9232;
        state = 128'h7f2c_3846_21c5_0400_a8a2_8710_2181_fbdb;

        #200;
        key = 128'h4694_7476_a337_e97f_b5bd_8048_0d4a_a5bf;
        state = 128'h4d86_6f66_88ff_4dc3_a7e3_60b0_52f3_d9e4;

        #200;
        key = 128'h4bec_1448_eb11_afe5_5575_f7c2_a070_88a7;
        state = 128'h0174_f779_e228_7292_2c17_0822_fe88_ecf9;

        #200;
        key = 128'hbd01_7462_b417_c43b_1125_9035_524f_cd7e;
        state = 128'h6e40_588f_a312_0324_0410_2f2a_c964_42c9;

        #200;
        key = 128'h0a55_479c_2b0a_47df_9a19_6a2e_b6e7_9618;
        state = 128'h2333_1e38_9d3f_59e3_ef64_f574_de6f_0041;

        #200;
        key = 128'he45f_fa31_b072_8f80_b2f5_99a0_993e_40e2;
        state = 128'h5267_97f8_a552_c2ab_3b2b_1468_bdb2_1a08;

        #200;
        key = 128'h054b_a033_05d5_4ea2_fd90_bbaa_b0c8_8394;
        state = 128'h2c02_1eb5_d116_53c9_d1ee_06fc_1c85_6377;

        #200;
        key = 128'ha8e0_dfd1_e764_84f4_643b_01c1_c05c_256b;
        state = 128'h1492_cde9_0ea6_3eb4_1acd_c956_4f2a_6bd7;

        #200;
        key = 128'h6a0b_07a4_c5b7_7d11_06b1_e30e_e208_6912;
        state = 128'ha5c0_1403_1d3b_4654_828e_55ec_9c18_786c;

        #200;
        key = 128'hb3dd_f797_b1bd_2407_e78c_6ccb_0c5c_11d5;
        state = 128'hac7e_17f1_b55b_4a53_83f3_9ec6_7646_6b8b;

        #200;
        key = 128'h8a4c_3c5d_10a3_f15a_7c69_11ad_3f1e_de9e;
        state = 128'h3a35_6714_3551_bebe_9746_1885_6763_0e10;

        #200;
        key = 128'hcf1c_0d77_5b8f_d1e5_6b0d_a596_7cc5_17c2;
        state = 128'heb4e_4c67_79de_cc8c_1a68_16e8_0d13_7a91;

        #200;
        key = 128'h7365_e822_7794_9020_73a9_b5f1_cd32_d75d;
        state = 128'hb6be_6c0f_a487_5d8d_42f1_96b5_5c74_dff8;

        #200;
        key = 128'h6c2d_4a0c_39a9_f6cb_7e84_7408_e150_5f8f;
        state = 128'h8d61_2a42_19b7_0e75_f400_438a_1c3a_679d;

        #200;
        key = 128'hc46e_f838_224d_f5e2_1bb7_4b37_a759_9bdf;
        state = 128'h0111_140c_b06c_f2dc_c8d7_f9e9_4600_34d2;

        #200;
        key = 128'hc3e4_2c25_81e1_e623_39d6_4548_40bb_ab6f;
        state = 128'hcc2d_3bf7_9a75_7a14_7abf_f697_cb15_09e6;

        #200;
        key = 128'h70e1_8673_983c_7b38_7ff6_c27e_6511_55eb;
        state = 128'hcfce_096c_9ecf_716b_59a3_3082_9fca_3f43;

        #200;
        key = 128'had50_98f1_5bf8_b54f_4735_6a65_e917_f686;
        state = 128'h4791_67f1_a03f_ce7f_df97_48ee_1c6b_349a;

        #200;
        key = 128'hf42d_ed60_ea3d_0559_97cb_86c7_4d21_f1e9;
        state = 128'h858c_4b81_a222_777e_2e20_ba70_2318_bc5e;

        #200;
        key = 128'hb001_b975_0afd_79e0_1dfa_acd8_e1a4_3fc3;
        state = 128'h44ba_9c43_815d_e49b_13f0_44be_56d1_1301;

        #200;
        key = 128'h4cbd_57ff_21cb_ab78_df85_51b3_bc6c_bac6;
        state = 128'h887b_3fd0_358c_b4b0_6f14_0892_d64a_1998;

        #200;
        key = 128'h58ca_e77a_8c21_a376_9721_b21d_5d54_cee7;
        state = 128'hea3a_632c_537e_c53d_d119_b7c0_7e72_3169;

        #200;
        key = 128'h9ce8_0af6_33ed_ba1b_87b5_4509_5ceb_08b8;
        state = 128'hd309_419c_0895_8052_15df_8a0e_806d_dc61;

        #200;
        key = 128'h1c6e_0bb6_b0fc_298a_e7fc_1a5d_e278_f8c5;
        state = 128'h473e_5774_9810_ed03_5fa6_5b7d_2bff_5b37;

        #200;
        key = 128'h6d41_c02b_e1c8_5cfa_9bee_3752_dc64_f768;
        state = 128'hfd63_5ec8_a044_4fff_37e4_34d2_9b51_cf89;

        #200;
        key = 128'h74cf_9ad3_0a0c_7855_8863_3d4e_f68b_4f2c;
        state = 128'h8eab_23da_50d1_042e_cfea_fd27_0eed_00e4;

        #200;
        key = 128'hdd7f_c6c3_a38a_684c_bac0_b9e7_c9c1_9c87;
        state = 128'hfbfc_a56b_1cf1_e2e5_87e2_eaf6_9d6a_9a64;

        #200;
        key = 128'hd15c_25f2_2cea_9e82_133c_359d_91b4_11a3;
        state = 128'ha0d8_9e68_6bd8_569b_e43b_2b4d_ccd2_653e;

        #200;
        key = 128'h0978_263d_4f12_3bda_902e_9a50_9ec5_a596;
        state = 128'h3637_4cc5_a380_9e94_a70c_6274_61fd_5800;

        #200;
        key = 128'h7c1d_1590_930a_5a53_930d_1a48_3ca9_638c;
        state = 128'h27a4_6071_8801_a30a_e08d_d9b1_b3a6_4dde;

        #200;
        key = 128'h3f84_2ab6_b27d_e766_c505_b468_23ea_3698;
        state = 128'h853b_bd3c_c2f8_50ec_8352_6272_885a_8f77;

        #200;
        key = 128'h8c1a_42bf_a6ed_81b2_0706_ec2a_929e_4c84;
        state = 128'h668b_7a50_285c_c290_ffc4_ebe8_a22b_b872;

        #200;
        key = 128'h5270_92b9_7305_00ee_2480_88c9_4daf_f2ea;
        state = 128'h19cd_44b2_e8f2_e494_a1ce_80cc_a28b_d1d7;

        #200;
        key = 128'hddf0_c98e_502e_cc1a_e983_deed_9bb8_ec0d;
        state = 128'h54e5_d54f_ac01_4080_db26_5ed2_4d09_9e44;

        #200;
        key = 128'hff66_3420_8eba_2820_6338_5bc7_058a_436b;
        state = 128'ha84c_6d92_5839_2ed0_858d_22e6_9338_4693;

        #200;
        key = 128'h7ccb_672c_03ce_cf08_5d00_9042_3247_36e3;
        state = 128'h37a7_aeb1_9b58_296b_5d5c_86ac_bfef_fd9f;

        #200;
        key = 128'h0dca_1f75_92ba_c3ab_1ca0_9d55_5085_1a6f;
        state = 128'h1cd4_fd3c_53e1_73b6_7e53_e86f_0e6c_372a;

        #200;
        key = 128'hd5a0_36f3_db02_acb6_c6ec_924a_5279_8e91;
        state = 128'hbf55_3e0a_8fb6_285c_3b61_c82c_56ea_8c2a;

        #200;
        key = 128'h4f2e_c874_726f_98ed_e825_5fdc_8fc1_e5b2;
        state = 128'h4cf5_1d8e_eb37_914a_7ad9_3455_26a8_0b29;

        #200;
        key = 128'h47f7_cdf9_8d52_32c9_e9a5_217a_e5f5_e21a;
        state = 128'h4dc4_3ad7_a015_3457_7a85_55b8_4315_3c3d;

        #200;
        key = 128'h5a12_a15a_60fa_ed4c_d43c_01ba_da27_e0cf;
        state = 128'hb383_1d8d_083f_f17e_af4c_4090_4645_8865;

        #200;
        key = 128'ha72e_0466_472e_496c_88cf_2ed1_11c4_b15a;
        state = 128'he647_b2c5_a47f_10a2_4433_694a_26b9_d405;

        #200;
        key = 128'h67ad_b644_0b16_4880_4e2f_12a9_cc05_28c6;
        state = 128'h3b53_6542_2de1_8dae_2de4_45a1_df5b_0999;

        #200;
        key = 128'hc832_d4c0_dbfd_8574_1a31_706e_fcd2_8d1e;
        state = 128'hadc8_e000_f671_8c2e_7f32_6613_8829_e006;

        #200;
        key = 128'hc31d_7cd8_ac2d_d733_fdd5_6574_604f_9f24;
        state = 128'hf35b_af31_2a69_2954_19a2_d67b_56bb_95f5;

        #200;
        key = 128'h6aba_7751_2280_d971_2593_f693_4ed8_2f2c;
        state = 128'hf4ea_c98d_6832_6221_75c0_9fff_793b_2cb7;

        #200;
        key = 128'hba5c_1135_e7bd_55e5_3836_4a51_3777_eced;
        state = 128'h0225_2783_0b4f_7afa_804b_10c5_17db_97e9;

        #200;
        key = 128'h4825_3327_030d_86f4_43b7_c28b_d3c2_ec33;
        state = 128'h93e6_f067_7238_3018_cc2f_fa0e_29d5_34b8;

        #200;
        key = 128'h921a_6cd0_18aa_c321_57f6_3f1e_e6ca_26ab;
        state = 128'h643f_3dca_26a5_4bfd_3629_e930_920d_fc25;

        #200;
        key = 128'h5f24_5dab_0aee_a081_b863_f62c_1839_6647;
        state = 128'hf985_0871_8204_1b01_6da4_d580_20f6_a6f8;

        #200;
        key = 128'h3418_79df_95e9_2add_9428_8edd_6ebf_1639;
        state = 128'h5566_c683_203e_3ede_3eaf_f1a1_910b_f2f9;

        #200;
        key = 128'h4961_41a9_bef4_5091_0024_64ca_ef5e_a383;
        state = 128'he196_8d0f_41cc_7a38_d2ae_b19a_a84c_36d8;

        #200;
        key = 128'h1148_a743_7d38_627c_8200_5d2a_cac7_2909;
        state = 128'h7d01_6c05_edc8_d410_330b_6ed2_c1d6_fdcf;

        #200;
        key = 128'h2490_5705_62e6_da67_00b3_5513_b796_0315;
        state = 128'h7016_b008_5690_7699_b170_2df0_dfe2_7ef7;

        #200;
        key = 128'ha955_b4c4_de7d_4dfb_3458_74dd_3516_790e;
        state = 128'he65e_95f1_7c88_015d_8e8e_182a_a53e_b48a;

        #200;
        key = 128'h2e2a_b77c_0f13_821b_3605_50ad_54e3_1124;
        state = 128'hfe6a_adeb_9237_a6ef_06a6_82f2_88b8_e699;

        #200;
        key = 128'h4911_be80_18c0_e58b_cd1b_496b_44db_9cdc;
        state = 128'h1c2f_54ae_de78_0d12_b9bf_d496_9ea2_a42f;

        #200;
        key = 128'hab0e_b023_c324_4bfa_6556_222d_a36f_faba;
        state = 128'hdbe0_ee7a_a1fc_f202_bd96_cf40_44fe_cc70;

        #200;
        key = 128'h629a_66de_002c_412e_6789_42fb_b14f_be6e;
        state = 128'h1a48_200e_f836_b5c1_65e8_76f3_6898_fd42;

        #200;
        key = 128'h0caf_2f0f_24db_e81c_7190_5990_80bc_d3fa;
        state = 128'h0cfe_af99_880b_0aa2_22a6_b373_e621_c191;

        #200;
        key = 128'hd255_36f0_813b_bd6f_e7fd_0fd9_0a27_54ce;
        state = 128'hc844_4234_7c88_6d12_ef7b_acc9_bc5e_6c7c;

        #200;
        key = 128'h79e8_0693_3b53_a008_6e90_5039_09de_20a2;
        state = 128'hf8df_143f_91de_64f6_9e90_ef23_4f98_660c;

        #200;
        key = 128'h92bd_a1b6_9229_dc77_f04b_a2d4_bdc7_f815;
        state = 128'h9849_30ef_57ea_8724_05fb_32b6_90dd_efbe;

        #200;
        key = 128'h53a8_8d4b_fb0a_29f1_b506_f10d_c8d9_eea9;
        state = 128'h4360_14f2_bbf1_e443_bc1b_53be_1c81_f156;

        #200;
        key = 128'h1c98_86e4_3869_f55f_81a2_5869_eb0e_0661;
        state = 128'ha265_e304_c4cd_24f5_d8f6_35d1_0508_7724;

        #200;
        key = 128'h95ba_3785_15f6_3467_41f9_2951_6a6f_66bf;
        state = 128'h219e_a63c_d44c_45e2_a83a_0b23_d6b6_cdb3;

        #200;
        key = 128'h4f44_6bb7_4c62_48c5_2a2b_3119_7882_633b;
        state = 128'h0a2c_f470_e881_cade_51ef_4d52_eacf_2796;

        #200;
        key = 128'h1fa4_3c87_31af_2f16_7a40_188f_2ae3_1bf3;
        state = 128'h983e_5c60_5c7f_4732_d78e_bd2f_b66c_12e6;

        #200;
        key = 128'he39b_0517_4327_8ba5_8b18_2e79_3ed1_bb95;
        state = 128'h575b_3561_262b_c9b6_67fc_3e46_83a2_c073;

        #200;
        key = 128'h0c36_52ac_859c_ee09_7c7c_c911_7a3b_4924;
        state = 128'h0712_68a2_846b_617e_8a4d_3179_a480_6e8b;

        #200;
        key = 128'hc5c4_a1d0_d181_6633_b304_9324_84a8_caa8;
        state = 128'h1bba_27f9_a8c2_7617_7300_a786_b3a7_0b0a;

        #200;
        key = 128'h7e3f_0e63_a153_e1f3_30c9_1b3c_5456_9ead;
        state = 128'h3876_3c07_cace_a467_4b95_af6d_dff3_dbd0;

        #200;
        key = 128'hc9d8_0096_95cc_9110_c1b5_2e44_aa27_83e6;
        state = 128'hea09_87a7_bc0e_28c0_919d_efac_f0e7_3a76;

        #200;
        key = 128'hb5a3_2b2e_c20e_ca01_be92_6a65_bdd6_4ce7;
        state = 128'hf707_5be4_0041_2379_08b5_72ea_7f0a_ecf9;

        #200;
        key = 128'hdc2d_e326_7c84_7a76_c07d_ab9b_31ca_d6db;
        state = 128'h958f_4d73_ca72_cd14_9e5d_a52b_bf21_b393;

        #200;
        key = 128'hd803_5ed5_cdb2_c89f_3ff2_aad6_0215_b55f;
        state = 128'h4f40_cc4e_1251_fd27_ca04_6264_40ca_6f28;

        #200;
        key = 128'h53ac_268c_904c_2dbd_0fae_e7f4_3202_0279;
        state = 128'h9536_4a5c_c8ad_9100_7b18_75d3_8b97_55af;

        #200;
        key = 128'h3ff2_eaf8_dc19_a37e_dbab_7429_a523_b1ab;
        state = 128'h5722_c28e_6406_6565_1202_4620_a7e0_4a73;

        #200;
        key = 128'h0664_04c6_64a9_f404_8495_5365_4843_1ad3;
        state = 128'h0f41_6289_131a_a809_cc40_b13c_4c5d_d31c;

        #200;
        key = 128'h9887_a569_5f82_0dff_95a9_ad4c_e79f_7276;
        state = 128'h4cbe_5196_173c_9620_df2f_79fe_d91c_6fb8;

        #200;
        key = 128'h3a11_17a4_775b_97a6_afa0_c876_88f0_72ff;
        state = 128'h27e2_514f_abc1_a093_fbe5_19db_175e_f24a;

        #200;
        key = 128'h8ec3_95bf_fc59_f4bc_59f4_ccb9_7dcd_8c0d;
        state = 128'h1f4a_f051_57f8_3888_06ec_5be6_f62e_1afe;

        #200;
        key = 128'h5d9b_a6cf_0142_2ecf_1468_409f_1100_1b97;
        state = 128'hcf1b_b19e_94b4_ed7d_c8dc_e78d_7d81_58d0;

        #200;
        key = 128'he3b2_4d0e_3623_8258_3691_4ebf_07a6_709c;
        state = 128'h05e4_a10e_1fca_763f_533e_cb5a_913a_331e;

        #200;
        key = 128'h3dcd_1166_5736_cebd_20fb_fe84_bcca_90c9;
        state = 128'h9b42_d022_d868_01d0_305d_b109_6b30_1338;

        #200;
        key = 128'hb04d_ea89_43ac_2c4c_4322_5820_8db0_31a6;
        state = 128'h0368_41e8_88e7_6976_63d1_b0e9_5312_195b;

        #200;
        key = 128'h4782_8a1b_36cf_1bd7_ca4c_22d5_ca66_5cf3;
        state = 128'h2faf_657a_9f99_509f_c83e_3944_ab5e_3789;

        #200;
        key = 128'h84b2_c655_0982_8392_78b3_e8fd_ceb8_b5cd;
        state = 128'he003_0008_4aae_f99e_54df_af6a_efa8_2c70;

        #200;
        key = 128'h6520_e70e_8ac5_9fbc_fdc5_3285_eff7_3131;
        state = 128'h7065_518e_f543_6754_ee19_5ef7_2be6_baaa;

        #200;
        key = 128'hde5c_74e0_7a5b_670b_19a3_c422_3e0f_a627;
        state = 128'h638f_9b9e_5b8a_b410_6d3e_cb2c_4917_d9d5;

        #200;
        key = 128'hde36_3b6a_3367_7d5c_b4ed_d916_cb51_8046;
        state = 128'h6f9a_7fdc_6105_78b9_816c_1f7e_7f79_7578;

        #200;
        key = 128'h36e7_0731_1a02_b46b_dcd9_283b_e664_ae0c;
        state = 128'h3c99_8dcd_bb12_f81f_d684_55d1_021e_79ea;

        #200;
        key = 128'h7415_c660_642c_1320_3f96_7c8c_0716_2607;
        state = 128'ha617_53aa_d7ce_7059_2848_514f_53ef_7ce2;

        #200;
        key = 128'ha52d_8dac_bdb7_77f1_5d65_6a7c_cde7_37d6;
        state = 128'h40c6_e922_d46a_3409_2eea_4dbf_89a9_be5b;

        #200;
        key = 128'h2b09_1724_9101_e1f3_3ad9_01a6_a13a_be38;
        state = 128'hae74_b7c9_2068_7c74_5624_50e0_96eb_c1dd;

        #200;
        key = 128'h9efb_9a3a_b2a8_edef_711c_e332_12dd_367e;
        state = 128'hcc7c_3b34_3f8c_6895_8363_02bf_ac7b_cd36;

        #200;
        key = 128'h06ce_42f2_df7e_7c6c_cae6_5e6d_1f28_d8b5;
        state = 128'hd641_8708_51d4_d3a1_cd30_6981_ae29_a811;

        #200;
        key = 128'h2362_693c_52ea_420d_4b0b_0132_6b87_73e9;
        state = 128'h19f1_62a8_57d2_aaef_ac3d_c3e9_a2e9_da81;

        #200;
        key = 128'hd2f4_bd84_6718_b2a9_29a7_f9ce_44d0_0b8d;
        state = 128'heb99_c9e2_53df_9205_4364_9b98_0769_39ad;

        #200;
        key = 128'h67b6_5f6e_5e55_81bf_34e4_3080_011b_223f;
        state = 128'hd6da_3a46_a7bf_cf0b_a46f_4476_6e0a_8031;

        #200;
        key = 128'h86ee_15a3_731f_521f_7af3_b448_b914_cf5b;
        state = 128'haaa6_f600_9a87_cefa_959b_9a39_6b7f_c585;

        #200;
        key = 128'hdf8c_0afd_8711_7be8_d254_74c9_8f5f_66fb;
        state = 128'h071c_2fb0_3ce5_c311_1e8e_e44c_2c26_23c8;

        #200;
        key = 128'h55b4_f7ad_d4b8_c3eb_fe1d_566e_6df6_8bc0;
        state = 128'h52eb_e613_5b9f_62bd_a153_14d7_d83e_c9a6;

        #200;
        key = 128'h03db_c21e_8830_c2b3_f19b_f7ff_c492_ce52;
        state = 128'he1c5_b422_ffb8_ed74_6e9e_859c_1458_6218;

        #200;
        key = 128'ha1b2_6c2f_3f92_8de6_6139_aff8_e64c_4a6b;
        state = 128'hbe0f_58ae_1a22_1d23_4ed5_2352_7e79_5daa;

        #200;
        key = 128'h5c9d_82c5_101f_b29a_32dd_c32b_df3f_afbe;
        state = 128'h86b5_99f7_572b_7860_5291_5cf0_e4ce_ebf9;

        #200;
        key = 128'h8880_8d29_48d4_5bc9_15ba_47d6_c420_08b7;
        state = 128'h5cb1_604d_6365_5c7b_0584_d0af_ac4c_b3da;

        #200;
        key = 128'h5e61_15ca_5ff3_d1d9_27d2_65e7_ca89_8181;
        state = 128'h8c87_53e9_625d_66d5_4ed5_8116_6da5_2295;

        #200;
        key = 128'h8d12_c1b6_a93b_8058_3566_d932_f05c_a023;
        state = 128'h783b_6e42_7292_4a59_ed05_e433_0e9a_c145;

        #200;
        key = 128'he76e_8eb7_dcac_d91a_8c23_ed44_1f35_786a;
        state = 128'hd44e_6041_d59c_6f9b_a60d_6902_76b2_1097;

        #200;
        key = 128'h4841_dd62_388d_6ff7_f45f_edea_3ec6_0c60;
        state = 128'h5334_f18e_ff74_8262_3676_d6be_be00_a11a;

        #200;
        key = 128'h65bb_a640_9355_aada_ef14_e760_d672_9785;
        state = 128'h0bc0_5d17_f273_9362_f719_7321_b28c_25b8;

        #200;
        key = 128'hf43d_b010_9586_0f81_24b9_7d1e_5bde_c78d;
        state = 128'ha8f0_c287_650e_f649_eda5_6be7_8298_e1d1;

        #200;
        key = 128'h3d1e_7d15_0f6d_425a_34d3_8b2d_3212_51f9;
        state = 128'h34fe_976f_cff5_4300_2ad5_ac00_6409_1e42;

        #200;
        key = 128'h1db9_0268_545f_b626_0fcc_e1f7_58ff_1ca3;
        state = 128'hf2c1_099b_7986_29d6_ae43_e56c_8927_5925;

        #200;
        key = 128'h68a4_d508_b1aa_4bf5_a231_1b40_ae94_d292;
        state = 128'h8a58_973a_b86a_a97f_ca0a_ad83_b4fb_55c4;

        #200;
        key = 128'hdf2c_c9c4_97be_d302_b701_ff09_36a8_c9a9;
        state = 128'ha8d6_8d23_adf6_c170_c7fd_1929_b688_ae9e;

        #200;
        key = 128'hb852_5ec6_3779_761a_a460_ed24_9e96_abd6;
        state = 128'h8e23_0b9a_8c9b_37ab_0c44_d953_1a52_0a16;

        #200;
        key = 128'h4470_61c2_f37f_d0a5_d403_bed4_e3bc_3f4d;
        state = 128'h5d02_445a_3060_c1f0_fda7_b698_a398_cf91;

        #200;
        key = 128'h3625_7cb5_7503_24ad_d2a7_c934_143d_3c83;
        state = 128'hbbb1_27f8_f03c_c240_d7f6_356b_4e14_9ac6;

        #200;
        key = 128'h8634_c4b5_9928_9df4_0fa2_d1a6_ae76_9baa;
        state = 128'h18e5_214e_ab50_81ed_a716_7b39_02f6_1925;

        #200;
        key = 128'h45b5_d83b_c6b8_de79_a9f3_03e1_4328_d89a;
        state = 128'h1e78_6b60_72ed_b77e_9fb1_4487_6969_9755;

        #200;
        key = 128'hb97b_dc2b_b5d4_b964_4a79_eb61_d5b5_f1ae;
        state = 128'h4fe0_c666_a9bf_8b4e_98a4_bccf_e767_b085;

        #200;
        key = 128'hbc8a_6bb0_83c0_2ca1_f843_cc39_003a_f254;
        state = 128'h6aa8_64a1_2344_ea46_f7f1_209a_7999_992c;

        #200;
        key = 128'h364e_8f6b_8942_78cc_f871_93d6_b533_19de;
        state = 128'hdb90_351d_b242_8077_983e_d20b_ebac_fda5;

        #200;
        key = 128'hbcc0_2a89_7c0e_e8fc_4d11_24ac_7dcd_d830;
        state = 128'h7166_272c_5083_a14e_9d2b_6669_c1e1_b920;

        #200;
        key = 128'hf6ac_2f57_7500_0af9_2eb4_f580_5d3c_ec9b;
        state = 128'h1f0d_f581_d9c5_bd56_553e_96a2_d2aa_c8e5;

        #200;
        key = 128'h06f6_18cc_3792_3224_bd1e_f4e4_d44e_ea40;
        state = 128'h270c_832a_f385_f5c5_1763_4cd9_761b_4235;

        #200;
        key = 128'hf8ad_71c7_b4f0_26fb_b9cf_20cf_711c_25f5;
        state = 128'h5822_8e83_9d95_2ba8_05bf_966c_ddb2_6000;

        #200;
        key = 128'ha026_4a50_499a_5a27_c7fd_3c55_22fe_034c;
        state = 128'h7b36_3723_23a0_2796_d0f6_4198_e478_70f3;

        #200;
        key = 128'hb686_61d4_46bf_01ce_290b_64d8_9e61_2b7b;
        state = 128'h0027_e15a_162a_fb9e_95fc_4b76_5e00_055f;

        #200;
        key = 128'h89ef_3b89_7ca8_9514_a2c4_2e84_0939_8c2e;
        state = 128'h8356_d248_8854_ef24_700a_0bd3_7147_79a3;

        #200;
        key = 128'h9f12_52ae_a3bc_54ae_f193_b940_2c72_bf9c;
        state = 128'h7e6b_2bba_98e6_d1c7_f4db_43c1_917e_d86c;

        #200;
        key = 128'h1cd1_ea33_1161_b52f_a8dc_afba_0d2d_71bd;
        state = 128'h102f_70e2_2a69_99fb_e130_e5a2_413e_2f2a;

        #200;
        key = 128'h8643_0ab8_e060_8bdd_8402_bca7_fae3_629d;
        state = 128'h66d8_5832_ad7b_625e_37fa_6b6b_b67a_ae26;

        #200;
        key = 128'h04d0_d014_07a0_07f8_5ec2_6e12_c017_e07a;
        state = 128'h939a_146c_b1fe_7210_7447_cb5c_57a5_ec0e;

        #200;
        key = 128'hff09_6cd1_309a_6aa1_a84b_a58e_2231_4f06;
        state = 128'h2138_a9f6_7232_305e_54a3_e6d5_8111_57ac;

        #200;
        key = 128'h63de_1494_7377_adb4_6722_871a_53f4_2fc6;
        state = 128'h41e1_95e6_a8ea_c899_9e94_acd1_ad1b_0a6b;

        #200;
        key = 128'hc122_5a5b_ccc5_5252_3e57_119e_aafc_7af7;
        state = 128'h47ad_3993_abd6_5523_d46a_8649_6056_82cb;

        #200;
        key = 128'he410_3f32_de8f_d17c_6a31_d8f3_d534_96fd;
        state = 128'hdd6e_6085_6cc5_1e70_84ca_3ad2_97a2_dbdd;

        #200;
        key = 128'h685e_1731_100b_695d_27c4_a3fe_99ef_46db;
        state = 128'h8804_3e1c_5a4b_b5af_d8ca_8550_a470_e25f;

        #200;
        key = 128'h64bb_42cb_7aa5_3c41_32e6_50d0_7b58_71fd;
        state = 128'he860_7a49_bca2_7624_6453_fe57_ae68_28fc;

        #200;
        key = 128'h3b65_4b57_1167_be45_d0d5_049f_8176_972b;
        state = 128'h1e43_1899_daf2_fb3f_5534_b98e_f819_6374;

        #200;
        key = 128'h93b8_c879_75c0_89e5_aeef_0166_e6d3_5931;
        state = 128'hb75a_bd8b_0043_76a0_2c7b_1144_4452_72c4;

        #200;
        key = 128'h171e_d26d_2f57_0dd5_0e4f_f0fe_4495_2416;
        state = 128'hced1_95c9_f02f_933c_e05a_a484_e60b_7f8a;

        #200;
        key = 128'ha7aa_782b_80e2_ffbd_0d02_4955_051c_9691;
        state = 128'h2567_c85a_791c_3737_bbd2_a24b_b9dd_f1ad;

        #200;
        key = 128'h0688_326b_c455_43d1_5b4d_d0d1_758c_25ca;
        state = 128'h4484_fa8b_5801_9d09_86b7_e716_b132_d914;

        #200;
        key = 128'h89aa_d4e5_562d_8378_a4e0_9ef1_8477_4b5f;
        state = 128'h3dfe_7cf8_bae3_d1c7_7d9f_e82e_eb3d_73b4;

        #200;
        key = 128'hf238_a69f_980c_443f_a87d_b5f4_1183_6b4e;
        state = 128'h7111_e48a_2b96_0671_fdf0_015e_c9a5_d814;

        #200;
        key = 128'h01ec_10d8_922f_f698_d288_058d_28e0_172c;
        state = 128'hb9be_4cde_1caf_f006_014f_815e_2baa_23f6;

        #200;
        key = 128'hceb2_50b5_021a_549a_caa4_ee66_ff27_d054;
        state = 128'h76bc_737a_11ba_72b5_c2c6_93db_3cf7_9414;

        #200;
        key = 128'hc505_eb96_5c7b_98e8_92bc_b44f_78c3_9be6;
        state = 128'h1973_1ac9_03b0_d122_b448_460a_8b87_e23a;

        #200;
        key = 128'h88e2_7b24_f807_0a67_3239_6f6f_486f_994d;
        state = 128'hba93_cdd7_78dd_1bbc_a720_0f1e_5a73_9908;

        #200;
        key = 128'h6387_11bd_8e1f_e927_a832_451e_21ad_4a92;
        state = 128'h28f1_8586_bac3_0b9f_0353_888a_26fb_eadf;

        #200;
        key = 128'hea8e_f77a_e19a_4ba0_72f4_8458_a051_0fc2;
        state = 128'hf424_0274_810a_ec52_052c_6af8_5c5c_5fc4;

        #200;
        key = 128'h8931_c1cc_9094_60ff_fb30_a71e_b316_a18a;
        state = 128'he41a_3cfc_c215_b7a9_a78b_93ac_bb97_ef0c;

        #200;
        key = 128'h6eca_9039_27c1_f744_af33_306a_af3a_2207;
        state = 128'h1e7c_7a2b_1323_f768_cebc_a5be_e73d_796b;

        #200;
        key = 128'h6509_9241_60b4_0e30_8902_1e5c_e2d9_754d;
        state = 128'he9e0_e7fc_9a1f_4107_02e4_aabf_23eb_5833;

        #200;
        key = 128'haff8_8070_c9ca_cafb_06e1_51ca_21f8_d18d;
        state = 128'h7fbf_85e7_22e5_edf8_dc58_3cc4_f4c1_8007;

        #200;
        key = 128'hc3ea_fe35_63f1_797a_08fc_5fdd_62bc_3f95;
        state = 128'h145d_b11f_48e5_dfe0_a0ba_5555_5976_8c4c;

        #200;
        key = 128'hf416_96f8_f2b9_4df2_b405_9689_b9c1_3ecb;
        state = 128'h21f7_e9d0_7025_40de_5911_b3c6_b5f1_1625;

        #200;
        key = 128'h2e21_7ef6_682f_343e_933e_0833_2b18_89ad;
        state = 128'hae45_5109_b751_ad7c_7475_3caa_304a_dce6;

        #200;
        key = 128'hf0cc_6339_6100_3ce6_7c91_7e12_787f_9915;
        state = 128'ha1c1_8dde_3b2f_3bef_aacb_3756_c1b7_38f8;

        #200;
        key = 128'h5c4d_5046_7fa1_0316_df18_b840_ac87_6df9;
        state = 128'h5334_92d6_ee15_a54f_1d61_31fb_cb29_aa4d;

        #200;
        key = 128'h1420_879e_20ac_2f38_ff54_92e3_92b8_2511;
        state = 128'hff8c_eaff_a1f7_a7f7_f4d6_9356_b2ba_5c46;

        #200;
        key = 128'ha659_2e33_e87e_48d8_b139_22e3_eecc_084f;
        state = 128'h2554_4969_f2c5_b6a5_63a4_53c5_b0fa_be29;

        #200;
        key = 128'h36a9_d7a5_9d31_6574_962e_ed75_d66e_3658;
        state = 128'h4ccd_e981_9971_fc59_a9e7_2c9c_9673_3400;

        #200;
        key = 128'hf2e5_5ea3_1157_14e7_83e6_93a4_2a48_261f;
        state = 128'hdd39_584f_5316_5420_1a10_a96c_da17_6736;

        #200;
        key = 128'h6b3c_f0d3_7a2c_ec51_faa3_7464_ce58_210e;
        state = 128'h654a_36b2_dfd4_b13a_02a9_cbf0_0093_a7d8;

        #200;
        key = 128'h4789_3d3b_442f_30e2_1bba_3cb5_f472_c434;
        state = 128'h55d7_b960_b96c_509e_1d0f_b64d_5f6a_442c;

        #200;
        key = 128'h7a48_5744_ad17_8c8a_5b43_45cb_1e2c_0bdc;
        state = 128'hac94_33b8_a9fe_4510_3d28_f885_526c_f5f7;

        #200;
        key = 128'hf095_8697_02a7_002d_549a_4b76_135f_dfa3;
        state = 128'h0ad6_8a2d_21a7_518e_a82e_9e53_78c1_2fa6;

        #200;
        key = 128'h950e_621e_6a21_4997_e38e_90cc_a3ba_ae6c;
        state = 128'hdafd_8fd0_6447_96ff_3748_0eb6_c935_ee8f;

        #200;
        key = 128'h1dec_1cec_0c61_5428_99a9_40ad_7194_d41b;
        state = 128'h4ebe_22de_065e_ae1b_7894_2d33_3256_7859;

        #200;
        key = 128'h524f_9d93_ab0d_6ae2_f1b7_6832_404c_bf9d;
        state = 128'h8d9a_3e65_b5c4_9e9f_b209_f42a_2efc_eb90;

        #200;
        key = 128'hb2eb_d005_3821_157f_81da_65ff_902d_fce6;
        state = 128'h94bd_00ac_2f85_ffed_fdfc_a9d5_5c0e_42eb;

        #200;
        key = 128'h7801_4c52_8d73_9b35_76b0_ca02_0d17_ea29;
        state = 128'h8dd2_7fa7_0754_87a3_738b_d173_c1d0_c50e;

        #200;
        key = 128'h94b7_1b8f_514f_01e7_4121_3cf9_7f72_934e;
        state = 128'h1111_5e0e_f00a_d861_3b1f_c162_4af5_d5a3;

        #200;
        key = 128'h8cc9_5e69_55fe_bbbe_cf60_57bd_ad84_95fb;
        state = 128'he7f2_f4e1_30a1_37ed_c6d8_27d8_85ca_6fd5;

        #200;
        key = 128'h8a38_14d1_2863_b442_30d9_7156_e077_48a4;
        state = 128'h8982_4ec9_4558_c7a9_918b_d1b6_953b_90e5;

        #200;
        key = 128'hf615_0da8_7306_7ca3_2c92_231a_57fa_45ff;
        state = 128'h7bae_f75a_8e08_a116_772c_2f76_c1a5_428b;

        #200;
        key = 128'hde2d_354e_a8c9_d9e8_d9ef_d957_69ca_149d;
        state = 128'h2f26_7fca_6885_a1bd_e403_92dd_15a4_fe41;

        #200;
        key = 128'h9026_e21b_e1e5_d5d0_d714_1a61_9569_a538;
        state = 128'h8041_1e11_1bbf_08b9_c045_515c_24f8_4c0c;

        #200;
        key = 128'hb7bb_20b8_243f_ec23_3b85_6022_f834_b85a;
        state = 128'h9c5d_fa38_2e75_0e87_ba6a_709f_c41f_0743;

        #200;
        key = 128'h2947_79ec_0175_5637_9c22_b80f_a96c_c36c;
        state = 128'h0057_b7db_2143_2519_ed18_0781_0327_43df;

        #200;
        key = 128'h590b_3cec_b5a5_9219_096e_e2cd_6926_9b0d;
        state = 128'hd0a1_eeda_e3dd_5926_6ad6_77e7_5d1a_9b70;

        #200;
        key = 128'h0951_b641_52bd_d73f_0321_8e6e_0a61_b465;
        state = 128'h9ebd_3941_e15f_54d4_46ed_df11_30bf_9700;

        #200;
        key = 128'h558e_396f_6894_4696_1292_d372_de09_a80d;
        state = 128'he026_eaa2_46fb_f4ac_fe18_9ac3_f824_dae3;

        #200;
        key = 128'hd164_1aa9_8b21_2d34_b5cf_2841_d681_2457;
        state = 128'hcc79_ab43_031e_441b_a887_ea17_1bdd_1fc8;

        #200;
        key = 128'h6722_df9e_da08_b7f1_74ee_dbeb_ffc2_b145;
        state = 128'h3b74_7a32_b7f2_2590_2b87_a5c5_c0d5_0a27;

        #200;
        key = 128'hb401_4f67_2f54_3776_0ca5_d101_f8e5_f7c9;
        state = 128'ha0a2_c476_9280_590e_e7fc_e6a7_efe1_957a;

        #200;
        key = 128'ha1c6_57a0_81e9_eb5d_a9b1_f7f5_3a59_a526;
        state = 128'h77ed_109c_3d41_8469_b3a5_8562_e2d5_49db;

        #200;
        key = 128'hf5c7_5c50_cd08_2c00_8431_28c4_fc50_fe7b;
        state = 128'h98ef_e7a0_6476_d37e_80b9_8d2e_5644_1998;

        #200;
        key = 128'hf3e6_e1e0_5fc6_7f61_0556_e269_2f45_d0eb;
        state = 128'h747b_d244_28bc_e7d0_60f3_0ab1_e13e_cd79;

        #200;
        key = 128'h4871_3aa7_d2cf_259c_89d4_5ca6_63c5_3a00;
        state = 128'h8f0b_331e_b57a_b2b0_fa1f_0e9b_520f_b5ff;

        #200;
        key = 128'h1804_6917_a051_6a0a_b107_9c99_14c7_431a;
        state = 128'h60e3_cfb3_80de_585a_b2c9_b9b3_bc97_9e47;

        #200;
        key = 128'hbe94_fea5_761c_d957_8de0_9683_ce58_703e;
        state = 128'h8654_10ae_ad6e_494c_0586_eb24_b5ab_ecc9;

        #200;
        key = 128'h7c6c_26ac_b076_b7a5_e6b6_01c9_fe94_783a;
        state = 128'hd584_5306_ce7f_ce74_3f4b_0920_440e_6738;

        #200;
        key = 128'h7339_1394_a2b6_2bad_1072_46e1_bd7d_efdf;
        state = 128'he438_affd_4d9b_2114_b6e9_4fc1_8392_2215;

        #200;
        key = 128'hb1af_c302_b9e7_7f80_0384_05b0_0f94_b334;
        state = 128'h18fe_402f_73f3_ed73_3cba_5b09_edda_c743;

        #200;
        key = 128'h5c40_2711_cfe8_e908_d56b_fb70_d6e8_b71d;
        state = 128'hcc6a_dba2_9084_8d4c_18c8_5afe_7690_6d43;

        #200;
        key = 128'h06de_73a4_4861_b898_d0e5_48be_c5aa_cb47;
        state = 128'hf592_3d86_f846_e3e0_b41d_5003_517d_1481;

        #200;
        key = 128'hac6f_e19e_08f9_d53f_b5c7_26e7_ae57_b9ad;
        state = 128'h2745_ff2d_f7d3_6081_b607_2c5b_4c62_cbe9;

        #200;
        key = 128'h98ba_f7da_49d3_f6cb_5559_9c8a_c377_8a07;
        state = 128'h346a_6f2e_b062_4044_3a7e_5f9f_9247_0b94;

        #200;
        key = 128'heaa8_e81e_bf20_01d2_845a_a13e_3d8a_53e1;
        state = 128'hf002_781d_86a9_92ff_d0e0_6f9b_b458_63ef;

        #200;
        key = 128'heb8c_cac4_d13b_ccb2_30a3_6971_0785_ee95;
        state = 128'h4b5b_c6a3_9ab0_a735_a3fb_db60_c006_4fa0;

        #200;
        key = 128'h53b0_a273_235a_4981_299e_7c3a_7f89_baa5;
        state = 128'hf855_8283_a634_80a8_514a_b7d5_c6a2_90be;

        #200;
        key = 128'h652f_911f_41d1_c0d9_8c48_4634_6a08_d599;
        state = 128'he10e_f861_13fc_1b6a_85db_cbbc_e6a7_a29d;

        #200;
        key = 128'hdf01_bba3_cadc_f6a5_d10e_24bb_de19_b259;
        state = 128'h967d_f53f_9b55_d960_6ba2_ca46_da4e_b3f1;

        #200;
        key = 128'h63f3_aedd_79d6_07d2_bf6e_8921_202e_a8a9;
        state = 128'h5f85_1d84_051c_4a0f_250d_d610_1005_9eda;

        #200;
        key = 128'h81a8_453d_a899_d0b3_a067_fca4_929f_5270;
        state = 128'h3a7c_3683_7d15_1d5b_1b57_cd9c_de22_e6b1;

        #200;
        key = 128'hcfb1_e5bb_7dcb_e33b_2e98_7e0e_a01d_6233;
        state = 128'h1401_de33_c579_309c_ab1f_97dd_69ce_8f83;

        #200;
        key = 128'hd263_dbb7_73ce_14bf_e4a7_7af7_d510_1ef2;
        state = 128'h520c_c8f5_81a4_5fef_1b0b_5f1e_23b8_24a5;

        #200;
        key = 128'h0b66_4970_e08f_61c4_dfdf_4d79_10e0_3cc1;
        state = 128'h7e46_89eb_72e1_f21b_5bb2_65cc_f17d_f5f4;

        #200;
        key = 128'hb96d_4ff4_7fa4_5858_f97d_9ef6_d5f9_456e;
        state = 128'h5b98_dc59_843a_2c14_c31f_de49_c5a4_ffef;

        #200;
        key = 128'he190_360a_6ff6_7df8_dc08_e844_a2f6_017d;
        state = 128'h70eb_e10f_53f6_5c2e_de2e_51b6_d55c_6d7d;

        #200;
        key = 128'hc741_3a37_5945_2bd4_74bb_1aa7_2332_2146;
        state = 128'h34e0_af45_c50b_2654_b942_6ea9_d3f5_3f5c;

        #200;
        key = 128'hb077_2c64_1e4c_1425_a88c_5137_60a9_76c3;
        state = 128'h75c7_3356_0b01_29d0_739b_c27e_7669_2cf8;

        #200;
        key = 128'h0e28_2c6d_6c5d_f8d8_b416_a081_83b7_4631;
        state = 128'h7dc4_5fcc_ec10_7248_48e0_3383_4b32_9c67;

        #200;
        key = 128'hc773_ad1c_2520_036b_361a_c0fb_6e96_656e;
        state = 128'hf555_c288_0e39_7e19_1efd_40e9_3003_ade8;

        #200;
        key = 128'hb6dc_02f9_d4a0_f771_91d4_8ab2_2f1d_d008;
        state = 128'h5ba4_eaea_5c63_a0d3_bd02_a161_ba56_d9f2;

        #200;
        key = 128'h8916_3d78_98a4_718c_f6bb_9c0b_bbb1_4dfa;
        state = 128'hc1a8_56bc_4248_bc9a_2287_41fd_894a_d1a1;

        #200;
        key = 128'hbcf3_40e6_cf76_92a5_e808_5ed1_19af_48c8;
        state = 128'hadef_e3f5_a049_b0f9_c46b_6cea_c6ad_3f24;

        #200;
        key = 128'h2965_4ed4_bbb5_e656_b017_3145_d565_9f85;
        state = 128'hd58c_5509_0db8_482c_a77a_eebf_e84f_6a81;

        #200;
        key = 128'hd6b6_8315_ca9f_facc_6433_3ba0_0644_1eed;
        state = 128'h904b_5506_641e_d98b_fe6b_b61b_04cf_d06f;

        #200;
        key = 128'hb620_e3e0_a43e_6ae8_8e70_233c_c64b_a536;
        state = 128'h2306_0103_997c_017d_e2b7_8da2_aea1_199c;

        #200;
        key = 128'h5f1c_5d9f_88e3_6317_de0d_888c_9023_9ddd;
        state = 128'ha214_2943_8daa_bb20_95ab_be21_54dd_6e80;

        #200;
        key = 128'h8c41_6475_9e1a_61d7_274e_383c_e0bf_cf03;
        state = 128'h1adc_fc61_9f7c_caa3_9e4c_d1ed_01ef_430e;

        #200;
        key = 128'h3895_ffdc_183e_6f2e_9759_43e9_b5fc_c55f;
        state = 128'hd9cb_ac0b_557e_4f0a_a2b8_4e13_733a_8570;

        #200;
        key = 128'h6005_f90b_ec09_2aac_6f06_c8d1_b68c_623a;
        state = 128'h0a4e_6096_51b1_ca3a_cd01_eacb_f635_af66;

        #200;
        key = 128'h9279_26fc_1053_0f9c_29c5_1ea5_98c1_e9c6;
        state = 128'h1dc4_c5bd_8524_47e0_1019_85c6_abc5_28d9;

        #200;
        key = 128'h4fb4_f0a7_2817_b3e9_d420_a2db_d384_b82a;
        state = 128'hd250_7a1b_bd32_dd5e_2401_151e_c1e5_f7bf;

        #200;
        key = 128'hedcb_f46d_2186_e102_940d_476f_3082_87a0;
        state = 128'h65aa_c935_a1ed_5ce1_8c89_1719_3c4e_87cc;

        #200;
        key = 128'habd2_35f1_d460_a585_4f4f_a499_627c_0550;
        state = 128'hec8a_4f4f_b7a2_5372_7359_44d5_63f9_9989;

        #200;
        key = 128'hf18b_8c1c_401c_7ec3_3aa2_debb_d77c_a485;
        state = 128'hbdec_658a_d7a6_923a_0c55_a24d_86ac_1952;

        #200;
        key = 128'h4d59_4df0_bbf3_30cb_24d8_eebf_0d61_4ed5;
        state = 128'hc23d_f39d_f555_565c_a608_3ac4_b6cf_f232;

        #200;
        key = 128'h7be0_17ac_4cd1_a649_3ade_4c8d_f3b2_7204;
        state = 128'hfff4_eef2_d70e_62f4_eaa1_da9c_5c94_e7b5;

        #200;
        key = 128'h4c81_96bb_1ba9_ea7c_542f_f9bc_8716_b655;
        state = 128'h4689_f48c_719e_3774_4c3b_89f4_9dac_47e1;

        #200;
        key = 128'h00bf_4360_0add_969f_23e7_42c6_163f_5bfa;
        state = 128'hc668_303d_e3a4_88bc_c2cb_10f1_2c2b_9420;

        #200;
        key = 128'h2680_73aa_8a7d_e716_f3d2_8dad_51ea_642f;
        state = 128'hd808_1c17_ebf6_fe6b_7000_f11e_2523_9cc4;

        #200;
        key = 128'h229a_9204_6287_41cb_eefa_69ba_e1c3_36c3;
        state = 128'h6d58_e715_18b7_652c_1b94_177b_f3e8_bab9;

        #200;
        key = 128'he08c_0c00_143a_00ec_0d41_2d4a_7056_1a4b;
        state = 128'h38c3_cec4_5592_2eb4_c468_5c15_02ac_80e5;

        #200;
        key = 128'hb45c_8ede_5b22_105f_2496_18d1_33d5_4fc1;
        state = 128'h1e11_e576_b4cc_922d_5b74_cf98_4614_962f;

        #200;
        key = 128'hb6b5_fbf7_d611_9739_69f4_7085_7ac5_3d2d;
        state = 128'hc8e3_030d_6572_2005_cdf1_25bf_4e3d_5b29;

        #200;
        key = 128'ha028_0242_a73c_0cb6_232a_909f_e1f3_cb15;
        state = 128'h7917_1466_2c4f_a68c_acd0_ebb6_129b_cb1e;

        #200;
        key = 128'h44a9_0dc8_de98_1287_a88f_af6c_7691_19ff;
        state = 128'he118_82c7_6f86_aebd_c716_555b_8f54_618b;

        #200;
        key = 128'h13e5_cbfe_ef2c_d99c_fa7d_cc74_03cf_cfa9;
        state = 128'hcb90_f4da_dc96_1751_e527_a8a8_8524_25c4;

        #200;
        key = 128'hec1e_61ef_8148_2ac2_4b0d_bb6d_c528_c843;
        state = 128'h6a56_417f_4050_102b_f0a6_cba3_75f9_c392;

        #200;
        key = 128'h7d76_0161_e226_957f_a784_5479_10a0_108b;
        state = 128'h5798_d0a1_52e4_116d_14f1_14e7_cfce_dd67;

        #200;
        key = 128'h10a4_4089_0be0_fc9b_f880_e1f2_5637_7e74;
        state = 128'hb5b8_8d90_ce25_3d9f_9581_ebc3_c158_4feb;

        #200;
        key = 128'hee8e_5900_ab3c_b2d6_393f_0c18_1f3e_65d6;
        state = 128'h79c2_871a_f7a9_3ef3_5f40_9a2e_1d99_c5e1;

        #200;
        key = 128'hcdd3_499f_2e7f_e2c2_f9fb_80a2_c2c4_a473;
        state = 128'hb6a9_3d7d_8df3_cc71_e65c_bea0_1d24_9e4e;

        #200;
        key = 128'h994f_dffe_d112_72a5_92df_32cc_0526_bc24;
        state = 128'hb53e_6684_11b1_a928_cca8_903f_ba72_a35f;

        #200;
        key = 128'h2808_b12b_4747_1248_98ba_b21d_1815_9893;
        state = 128'hea46_93d4_741a_e861_2b94_f8ab_c86f_05cb;

        #200;
        key = 128'h01a3_9adb_d3e2_e02b_b15f_34eb_ea7d_ceda;
        state = 128'h61fd_1c76_1cdb_1af4_6aa9_7568_7508_65f4;

        #200;
        key = 128'h3928_2824_6448_c6c0_617f_9ee7_7f8f_ba61;
        state = 128'he7db_8902_2169_23fe_bb31_b07f_e770_2725;

        #200;
        key = 128'hddca_9117_9b5d_cd51_3be8_cf9d_7591_6a4e;
        state = 128'h42ca_d875_e278_6cc9_7121_e546_6c6a_81f8;

        #200;
        key = 128'hd2f8_3520_8b80_dcac_d5de_f081_5ac8_c6c7;
        state = 128'h83d3_91f7_9536_65a2_249e_f8d7_7024_daba;

        #200;
        key = 128'hbe50_8723_4775_1d3b_debc_a0d3_3415_ab38;
        state = 128'h8c30_bf51_9cc7_d2e1_8ee2_00da_2bd5_965b;

        #200;
        key = 128'hac6b_9849_fbbe_8232_efac_a0e8_a967_3fd3;
        state = 128'h0636_2892_8020_f8cd_3c98_8fd4_9d38_eb12;

        #200;
        key = 128'h68d1_c1d7_b9df_a908_1b5d_1465_3ae9_ea9c;
        state = 128'h3989_337e_62e9_375e_6ac7_50fa_85de_a929;

        #200;
        key = 128'hf1e1_fe22_5693_5b3b_3738_a780_17cd_8837;
        state = 128'h0cab_9627_4492_427d_830b_977a_4ef8_9067;

        #200;
        key = 128'h61fc_1717_1914_684a_e883_f628_0983_939a;
        state = 128'he056_edfd_78a9_f0c6_61f2_745f_1ba6_70c1;

        #200;
        key = 128'ha703_f65f_f625_6751_d003_0b40_a797_4bdf;
        state = 128'hfb21_19e7_8b9e_0fa2_1b5e_be3f_79f8_5596;

        #200;
        key = 128'h9865_7a65_0ee2_57bb_21dd_b681_c231_bcec;
        state = 128'h67d3_57d1_6045_f1ba_3acd_dd43_794d_59c5;

        #200;
        key = 128'h02ea_ba4c_b9ed_0d7b_47f0_51de_7551_42d2;
        state = 128'ha3f9_4937_9b13_57d2_9fbd_4e8e_f1b4_a70b;

        #200;
        key = 128'ha3f8_4d65_0b73_1eb8_d47a_a40b_4006_18c1;
        state = 128'h637a_88af_6793_3550_c6b0_eb7a_339b_337b;

        #200;
        key = 128'h9812_ecb5_61a7_b359_133a_53f6_a417_de8d;
        state = 128'h3e52_d0f1_c7c8_b6b9_4d63_4ad6_a341_f06f;

        #200;
        key = 128'h0ac2_5735_3168_ac0b_cab4_d73e_0a89_67e6;
        state = 128'hf436_cf09_de8b_db98_c5e7_4217_a5b7_06e0;

        #200;
        key = 128'h2fa2_0e21_a317_3711_3d16_3778_de1e_4977;
        state = 128'hbcb6_facc_d601_331d_13e8_48c8_6036_2a6e;

        #200;
        key = 128'h39fa_3820_d27d_3bea_d453_80e0_543c_b45c;
        state = 128'h8f8f_6bc6_925d_c70e_f9c2_a7f6_ab6a_39f1;

        #200;
        key = 128'hef23_39e8_e92e_23c7_3fed_34ac_589b_fc19;
        state = 128'hc738_b258_9d89_6da0_393d_36d5_9059_3daa;

        #200;
        key = 128'hec27_75a5_9726_f979_bbcc_d3be_0d07_9e65;
        state = 128'hc332_552b_971a_e3ff_7fff_5f7d_9124_6497;

        #200;
        key = 128'ha426_fb5b_cc49_88a0_31a8_e695_56a5_8213;
        state = 128'hb7bb_9a3b_b0fa_b019_f51a_7461_8388_5fbe;

        #200;
        key = 128'h93a5_ea07_0af8_ffd1_c0a5_4501_9bc5_0162;
        state = 128'h50ca_7d2e_c5d4_8f9a_6957_02b0_00a5_5a2e;

        #200;
        key = 128'hc2ec_b8cd_955d_9040_5d72_a624_489f_4880;
        state = 128'hc346_6b41_ed2d_6807_a39f_6a68_8c95_ace3;

        #200;
        key = 128'h5b0c_d7de_ad51_5143_f8df_524e_5e96_8594;
        state = 128'hbb37_4af4_b0b7_9d95_defe_2cbe_c869_2dda;

        #200;
        key = 128'h45d3_ffa9_0189_704d_e0b4_7a04_8972_e466;
        state = 128'h1ad5_3950_5987_1dee_9914_71ce_7649_8d8c;

        #200;
        key = 128'h536c_153a_fd13_0e61_8503_fc9c_6fa6_b3be;
        state = 128'h5fa6_fa10_fd62_7b9a_d579_3892_7020_4889;

        #200;
        key = 128'h0ca7_f801_a3a6_de26_24df_4083_63f4_fda9;
        state = 128'ha7dc_5db2_5d21_2785_9e30_cbb3_fa4e_ac24;

        #200;
        key = 128'h3fcf_eceb_e651_4181_0aca_5152_28f4_d2a9;
        state = 128'h4c04_a22b_5ab4_48bf_fac1_8356_ff01_ff15;

        #200;
        key = 128'hd822_7ac8_a0e0_803e_d1ca_6d3d_83cf_25d8;
        state = 128'h06d1_734e_dd8f_a99b_2cad_eb8a_ded0_be59;

        #200;
        key = 128'h9902_d5ea_c0aa_728c_825f_a811_8f07_70b6;
        state = 128'h0076_935e_f3cf_82ff_e58a_91c0_123c_6870;

        #200;
        key = 128'hae51_5767_f17e_d87a_ad2c_5bdf_e466_2895;
        state = 128'h841d_18eb_8e8c_cba0_d90e_8cb7_b07b_88ad;

        #200;
        key = 128'h7a4a_30ac_6916_3f33_7a45_f2a1_6db2_83a0;
        state = 128'h0c37_1618_a2e6_d29f_c4b8_840a_9f5d_ba51;

        #200;
        key = 128'h8623_5deb_d95b_0ebc_6d93_3d76_b10c_9fa2;
        state = 128'hb1a8_a159_8083_3ff3_22e9_3904_c032_a0fc;

        #200;
        key = 128'h25e7_3b75_cc27_7e09_b413_1e98_8b2c_549a;
        state = 128'hbb58_d663_fe3f_3afe_d5a3_ce9d_0902_15ce;

        #200;
        key = 128'haab5_d4df_748b_67dd_df96_8c1b_5958_8ce6;
        state = 128'h40a3_afd3_7efc_f56d_34a3_8a1c_147e_2839;

        #200;
        key = 128'h4335_4925_a8ab_d220_1dbe_6eeb_b7fa_5ec6;
        state = 128'hba50_f4a4_c051_db85_f1ea_f740_75ee_42d0;

        #200;
        key = 128'h5e8f_51dc_40f9_887b_63fd_8414_9c57_4b15;
        state = 128'ha605_574a_7154_1cdd_d21c_13f5_ef32_3c30;

        #200;
        key = 128'hb6f6_ecaa_8f6a_18e4_654a_d65f_530c_b774;
        state = 128'h99e4_b927_4616_86fb_9be0_bba3_a9eb_5dce;

        #200;
        key = 128'h7dfe_98f6_26e2_7b25_dc4b_9923_cd48_7a5b;
        state = 128'h86c7_3e0d_e4c9_c7b8_8ecb_e106_0d66_f3c0;

        #200;
        key = 128'h2341_f83c_0a4c_f2bb_c323_d90e_945c_d5ad;
        state = 128'hacb9_2c89_577d_e796_dc3b_2d25_9c37_e410;

        #200;
        key = 128'h59bb_d529_4a1b_ecac_0065_d0a1_f848_3d33;
        state = 128'h077d_50d6_1f3f_543b_040e_f41c_67a3_099a;

        #200;
        key = 128'he68e_4bef_d7c1_361b_cb12_07fc_5676_fc58;
        state = 128'h2308_5fdb_a1a5_c5ea_3da2_bb42_3e85_90e0;

        #200;
        key = 128'hc253_d0f8_b94b_4b98_0879_ecbe_9bc0_7655;
        state = 128'ha05e_e99e_6054_8f8e_5ae0_be41_0328_a3ea;

        #200;
        key = 128'ha23b_847c_1681_9b42_8362_886a_c577_4075;
        state = 128'h2ae6_b7e7_870d_41c8_4e82_3877_f4c9_2272;

        #200;
        key = 128'ha523_bf46_f1ce_1877_bc2e_bb89_f23a_6a5e;
        state = 128'h3e6b_b7bc_92d7_a774_d36a_d02a_1d0d_4610;

        #200;
        key = 128'h54eb_d64f_7a6c_913a_4539_094b_7af4_f2b9;
        state = 128'h4def_eae0_9117_f0fe_605e_8661_be92_a946;

        #200;
        key = 128'h08b7_34fb_d548_3e91_39e8_bbe9_002d_93c4;
        state = 128'h60ab_b214_147a_8ba3_c9b2_a8f1_3c5f_91d3;

        #200;
        key = 128'h0809_2d3a_5bc0_33a1_23c6_a4fe_66b8_ef8d;
        state = 128'hb92d_4cbc_58c5_ea48_c0f2_7c71_733b_aa18;

        #200;
        key = 128'h42e5_c7ce_366a_416b_5d7c_0467_894b_4e83;
        state = 128'h56ca_3fe8_c215_b04b_af5a_faf5_7ebe_3c53;

        #200;
        key = 128'h264c_278f_7aa4_e55b_a056_b1b7_3953_d40d;
        state = 128'he82e_160b_81fb_c984_b2e0_05d0_7f56_b408;

        #200;
        key = 128'h6b60_0996_9cbf_0579_310b_8f05_72a6_fccd;
        state = 128'h7b24_215d_9dd8_4945_c2b4_a36d_004b_87b9;

        #200;
        key = 128'h64cf_fd9e_738d_907a_01cd_e8a1_c1f1_382e;
        state = 128'h35b2_673b_954f_8a3f_d00e_5323_16c2_aae6;

        #200;
        key = 128'hd3fd_ae63_8b4b_e3ca_56cb_2dff_011e_355e;
        state = 128'h7067_5701_e677_7f36_6937_9ec4_33fb_da31;

        #200;
        key = 128'h488a_df6d_c2c3_3ddc_2e2a_905f_1499_c3ab;
        state = 128'hfd65_27aa_42d3_f116_ba3a_9794_a7ae_182c;

        #200;
        key = 128'hf737_741f_c464_9560_e80a_ff5e_ccfb_b749;
        state = 128'hc6bb_2620_79e2_c232_f5aa_3ac9_4a21_72ca;

        #200;
        key = 128'h3ae7_c0dc_9d86_9a55_c54b_a6c6_3187_7ab9;
        state = 128'hfae9_8712_41d6_e756_5709_f40e_de9c_e5de;

        #200;
        key = 128'hef4b_1803_804b_9911_332a_a153_2af7_c4c4;
        state = 128'he57a_2bb7_c8f0_54bf_a588_45c7_d3b8_3e97;

        #200;
        key = 128'hf065_8236_c808_023d_8fb7_55cb_1605_cbff;
        state = 128'h2282_02f9_40c1_9bfa_d27a_3fff_1fae_98d0;

        #200;
        key = 128'h03ff_7482_3fc1_9ab9_6e72_ca91_6834_cb47;
        state = 128'h12d4_3d8a_0b15_96cc_02ad_07ed_853b_968f;

        #200;
        key = 128'h0a2b_be0d_ba04_92c9_b18e_27ce_1e31_8f9f;
        state = 128'hd49d_b444_b16d_d11e_914d_24e4_b6a9_0887;

        #200;
        key = 128'h87b3_225a_5343_9fba_2d90_fe59_9187_4678;
        state = 128'hb540_c40f_6be2_f67a_ab21_cd78_2557_3104;

        #200;
        key = 128'h92d8_5173_838b_4e4d_1659_8585_42a1_4d92;
        state = 128'h6ea0_3250_7962_ef7f_292f_1be6_96df_a635;

        #200;
        key = 128'hc169_c438_f5bb_19cb_827f_67ba_20e0_da3e;
        state = 128'hca39_5d25_ea0b_20f5_04cd_36f6_319a_5498;

        #200;
        key = 128'habaa_f310_6133_ad1d_4a45_ab7e_b30c_c4e9;
        state = 128'hcf23_e529_a00b_cbd8_1a2a_28d4_488f_63ad;

        #200;
        key = 128'h5954_2bc1_465b_294c_686f_aeb7_1e1a_7147;
        state = 128'ha4d1_5f84_c830_0b76_fcf9_0185_ba39_ef8f;

        #200;
        key = 128'h29b2_8b71_0541_7d4c_58a7_137a_abe5_f9d6;
        state = 128'h0f64_1fc1_43a9_a3fa_baed_0f41_8cb0_99dd;

        #200;
        key = 128'h6857_ced3_ddf8_07b7_c5ef_41b6_7042_4e89;
        state = 128'hebf1_cdb2_7963_b7f8_6df5_ffb7_9917_f64f;

        #200;
        key = 128'hf685_283a_053f_62d8_7e5d_fb06_1583_2087;
        state = 128'hf1e1_b3d2_fde5_5a32_5057_762b_e68c_ca07;

        #200;
        key = 128'h7501_8f98_263c_300b_84eb_7ff4_7726_014b;
        state = 128'h4645_68d7_f500_2fc0_9a92_2c55_16c1_98aa;

        #200;
        key = 128'h72f6_304f_8568_bb69_c0c9_4f61_751f_2753;
        state = 128'h7d83_f9e7_16e5_321d_d2f2_faf6_ce78_e5e9;

        #200;
        key = 128'h9548_6466_69ba_3e41_2bdf_4f65_7211_de89;
        state = 128'h79fe_9b3e_4e53_2445_150b_d8e9_1008_2fea;

        #200;
        key = 128'h0a3d_2517_d2f5_b4de_86af_b739_64a8_8d11;
        state = 128'h44ba_7e8b_6429_b49b_16f5_b618_b17d_6dfe;

        #200;
        key = 128'h7a2c_3b09_94a5_f800_df35_6e53_9d02_8204;
        state = 128'h9ee6_2a82_cc33_e7e7_d317_c456_29bf_742e;

        #200;
        key = 128'h6d8e_4860_d322_88db_6ac8_652f_6edd_3f71;
        state = 128'hfe08_928d_0970_b0f8_c5bd_737b_4642_1050;

        #200;
        key = 128'h6ec2_701d_b7e5_563a_230e_2a85_da89_ca8a;
        state = 128'h9775_d18a_32fc_0684_c1c5_30df_eb04_d380;

        #200;
        key = 128'heefd_cf4a_5418_7d5a_05d6_fc93_52af_613d;
        state = 128'h4317_6d5b_9553_1d1c_b4b8_3957_cd43_b274;

        #200;
        key = 128'h4eeb_84c1_4881_c9e3_64f5_c9e1_772a_a50d;
        state = 128'h7460_f441_706d_d6a2_85c2_aee7_4df8_7ca8;

        #200;
        key = 128'h5b3e_7fa1_cdf6_375f_f977_2269_9163_1427;
        state = 128'h5de2_c244_e1e5_4a7e_11c6_084c_f0a7_5ee8;

        #200;
        key = 128'hae6a_aabd_b4e1_fbdc_5571_4ea5_15fb_a7c9;
        state = 128'h9052_d0ee_cdb0_346c_c231_3c94_ea43_6478;

        #200;
        key = 128'ha94e_09bb_d69c_77f9_186a_84c6_a00c_dad9;
        state = 128'h6436_b5d7_3977_83df_d14b_ae64_affd_7478;

        #200;
        key = 128'h71d3_37de_5298_1bdf_11bd_9666_8bdc_200d;
        state = 128'h0c7c_8095_11c5_6b44_038d_d878_a9fd_33af;

        #200;
        key = 128'hff6b_05d9_279e_a140_9991_9802_0ed8_d25f;
        state = 128'hceb1_dd9f_a900_e9bd_03be_3ddf_f4e0_81f0;

        #200;
        key = 128'hb008_78d1_5faf_8e1f_8a8d_5a24_dff0_bdce;
        state = 128'hb53d_57d4_411a_aed7_de0f_e3b0_afb0_28cf;

        #200;
        key = 128'h238d_efb6_35bb_882e_e18b_cd39_645e_b789;
        state = 128'hcfed_82f1_62f1_96fd_c59f_83fe_e95b_574e;

        #200;
        key = 128'h5fa2_5f61_e64a_f7b2_eff7_33ed_df4c_e77e;
        state = 128'hcef4_c6b6_833a_1340_e9a9_dbe8_ce9a_8d9d;

        #200;
        key = 128'h1b7b_4b5b_9063_4964_babc_246d_3a7e_3e35;
        state = 128'h20cf_3115_713c_5769_9017_42e2_0934_1688;

        #200;
        key = 128'h38a6_2d50_be2f_7643_336d_8b0b_9e23_2598;
        state = 128'hcc73_482e_0776_b127_f69f_bbd8_4242_4e65;

        #200;
        key = 128'h2cd1_f686_8392_e32d_a761_d8f1_43a7_6120;
        state = 128'hf66f_c357_2d76_e09f_5aa1_bb61_770e_faf6;

        #200;
        key = 128'h5540_449f_0f92_57c3_62c9_d1d9_951a_0d4a;
        state = 128'hc546_bf4a_c07f_2ee9_e764_adfd_c7d9_8ca5;

        #200;
        key = 128'hdf97_03ca_2b40_2c6c_0514_3ac1_04ad_88e9;
        state = 128'hb8ec_82d3_a184_436a_5801_da39_f6e9_44d2;

        #200;
        key = 128'h61d4_8dde_6745_f1cd_850b_67e9_ca00_5d8b;
        state = 128'h020c_dc8a_43cb_6ebd_b535_d969_f11b_0a15;

        #200;
        key = 128'h4cfb_fcfe_01e0_477e_4ef1_bf89_b7db_5705;
        state = 128'he6e6_cdc5_e9a0_66e4_5a14_a46f_c50e_83a4;

        #200;
        key = 128'haa66_3167_b64e_5ef6_9440_802d_a97e_05d8;
        state = 128'h914d_d27d_de8a_948c_ba29_f3e7_f08e_f8f1;

        #200;
        key = 128'h95bb_0200_99b5_a449_047d_d158_7b9b_ffd1;
        state = 128'h4f4d_0495_1bff_7627_ed0d_2adf_8efa_55cf;

        #200;
        key = 128'h2000_b725_3d7c_a41d_c898_a5b1_1b34_1669;
        state = 128'hcf77_2933_f799_1165_f68a_4ff1_37c3_04a3;

        #200;
        key = 128'h9f32_efb4_e735_61f1_cec3_afe9_8009_671c;
        state = 128'hbf16_fadb_cda8_493e_adf9_ba83_3ca5_b92b;

        #200;
        key = 128'hbf07_99ad_cfe2_3dc7_40f5_9fb6_7f5b_e26a;
        state = 128'hf081_8602_71f4_2194_5ad1_2681_8ec3_201b;

        #200;
        key = 128'ha0ab_5120_7d01_b5da_45d7_60c1_218c_fc04;
        state = 128'h0ab0_b4af_203f_5eea_2132_795e_a6cf_be00;

        #200;
        key = 128'h635f_5902_3237_cf14_f7a4_25c0_c4d9_e994;
        state = 128'h85ef_bd88_42ff_b260_504b_11b5_a4ab_ce91;

        #200;
        key = 128'ha615_3edd_c6a2_6de5_51d2_eef0_c1c9_6cec;
        state = 128'h467d_7db8_0594_40d4_d575_9627_d488_2936;

        #200;
        key = 128'h466a_9121_77bd_1436_7147_3e38_75ff_21e2;
        state = 128'ha00e_bfea_0433_0fa2_e89b_d36b_aefc_e4f8;

        #200;
        key = 128'hd4c1_d79f_0299_91f9_3113_a420_6d96_99fa;
        state = 128'h1281_604e_a1cb_bc4b_b4e7_f3c3_f646_8cb1;

        #200;
        key = 128'hbe83_60b0_338d_26bb_d663_a2cb_ba47_b0de;
        state = 128'h605a_f905_4df4_bd7c_0234_e9f3_fdec_74c6;

        #200;
        key = 128'h436d_485e_118d_f044_0576_5768_fcc2_4de8;
        state = 128'ha390_f3ec_6d3f_e02b_902a_6a39_3969_eb0e;

        #200;
        key = 128'h82e4_b305_9168_3e2f_2ede_22d1_77c8_eeb2;
        state = 128'h35fb_e584_f69d_5f2e_5373_f046_0d89_8a6c;

        #200;
        key = 128'h6fb7_7359_c5d2_54af_478a_a181_0609_205a;
        state = 128'he000_809d_bfcc_e60a_9c6e_6845_c24e_2fd7;

        #200;
        key = 128'h45c7_45ee_4c94_27f0_0886_ddeb_1bed_8857;
        state = 128'h1312_be78_61e3_f1c3_713e_3ca8_80d6_8697;

        #200;
        key = 128'h734b_d1de_a082_f0b7_4e11_9307_8a2e_29cb;
        state = 128'h5578_8952_332c_98f3_eb82_c057_407c_2cc7;

        #200;
        key = 128'h7fa7_32f5_d452_fd0a_248e_54c1_5d80_f543;
        state = 128'hdf3d_de5f_9e61_8d95_6d9e_229a_954b_7946;

        #200;
        key = 128'hc9f6_36a4_5471_c1ee_bb28_5a7b_a113_b62a;
        state = 128'hebf1_8864_d69d_0736_39c0_ff11_d5f9_d83d;

        #200;
        key = 128'h5a32_164f_c4b2_cae9_5a89_1d31_edce_98ff;
        state = 128'ha22b_d7a3_e873_cf76_e085_d52d_1af9_f5be;

        #200;
        key = 128'h1866_1cb5_a759_d821_a893_95d1_fc69_2c96;
        state = 128'h7fac_430c_a4e6_2232_613d_f53a_a9e5_51e2;

        #200;
        key = 128'h056e_60ef_9fce_97fc_fb3d_4f20_cf8e_7446;
        state = 128'h8f1d_bd0a_0f72_5bb6_3749_8a19_1771_3676;

        #200;
        key = 128'hbfb6_5ab0_c930_6c6a_0811_31e6_4f24_c70d;
        state = 128'h5477_743c_43a1_24dd_6437_5ccb_b1cd_e8dc;

        #200;
        key = 128'h4fc4_3b03_0204_14c4_4297_bb80_4e5b_54e9;
        state = 128'h9bfb_c4a3_5cfb_7596_4693_888f_a99c_baef;

        #200;
        key = 128'hdcbf_4880_79f3_fba5_cd45_48bf_2b81_8619;
        state = 128'h5e84_1165_f28b_40bc_3e3d_6f72_0c9f_274e;

        #200;
        key = 128'ha942_9681_4235_ce8c_84f5_11f7_7fbf_7563;
        state = 128'h68b1_347a_1282_b835_a300_02c8_50ef_156b;

        #200;
        key = 128'hb8fe_579c_33a9_301a_99ed_8078_0a92_0c5d;
        state = 128'h9e66_bc14_6f43_2cb9_08d9_660d_e4bb_889b;

        #200;
        key = 128'h80b5_3fde_9be2_849e_5752_5d7f_af66_9917;
        state = 128'h38fd_16fb_5b79_7e25_56c4_85df_7408_76db;

        #200;
        key = 128'he00d_4db2_ce4e_8ad4_f816_099e_356b_52a1;
        state = 128'h3618_7f0b_377c_7312_219c_1136_18fd_ec0a;

        #200;
        key = 128'h4c1e_fa2a_d796_e3d6_f24b_2960_b532_2f05;
        state = 128'h4034_f4a8_c175_aea9_6d23_1c6c_4800_1887;

        #200;
        key = 128'hb92e_2a56_7723_8e9d_fb72_1080_2ceb_0353;
        state = 128'h7712_ebb1_bed6_0119_2a44_ee3a_6be8_4dea;

        #200;
        key = 128'h567d_790d_6a38_a1f9_50ae_2d80_268b_549f;
        state = 128'h1a25_2b0e_4ffd_41c2_9af4_fb2e_c0e1_1780;

        #200;
        key = 128'hde45_7a26_26b7_55db_03b7_99aa_0d6b_9735;
        state = 128'h7125_4de6_9695_f5b3_59c5_31a4_ff49_4981;

        #200;
        key = 128'hdfac_ee31_13f4_699d_88ed_08f9_d38d_f2b9;
        state = 128'h3d06_db17_bce1_5806_6d5a_7e88_2f65_fafc;

        #200;
        key = 128'h9281_05f8_43b3_3303_69ab_7b74_8283_367f;
        state = 128'h55b5_af1f_bc8d_b822_a482_2e51_2da3_6977;

        #200;
        key = 128'he798_f2b6_7d82_a445_4cd1_30fa_51c0_d093;
        state = 128'h7e52_b9a7_edb5_6220_3f5e_abf2_a03f_a05c;

        #200;
        key = 128'h36e2_e898_0f54_6dc3_c32c_2f29_475c_4b66;
        state = 128'h6dae_b5f5_56a8_9c6e_3d7c_9144_ee02_1193;

        #200;
        key = 128'h2951_8cf4_6a2c_b628_8a3e_db5f_fea9_b9bd;
        state = 128'hb26e_60a0_d885_44c9_4bb9_4623_5bad_7feb;

        #200;
        key = 128'h9ffd_7a8f_8ea5_8ba1_d35d_fd7a_81cd_acad;
        state = 128'h1e87_a64a_98ad_af04_c7d7_0ea4_e70b_ee18;

        #200;
        key = 128'h3e2f_d58c_6f79_1eb5_c061_b064_0f70_e80c;
        state = 128'hbacf_6689_5b7f_6f62_e191_bcd2_ad0d_cad6;

        #200;
        key = 128'h82ad_1fc6_bd9c_0970_5928_75e7_649d_c444;
        state = 128'hcf68_133b_4442_4735_c981_1485_72eb_ab0b;

        #200;
        key = 128'h6795_4d91_4259_a124_52b7_ebf2_8552_fc18;
        state = 128'h6b67_8659_3a82_b6bb_dc57_1b77_62b3_2cb5;

        #200;
        key = 128'hb5db_178e_6ab5_e206_7791_5f15_1324_9fa0;
        state = 128'h9042_f8e8_d627_8e3d_f961_08e6_61ab_808c;

        #200;
        key = 128'h8b39_3b20_5375_f7a1_d6d5_fd46_35ab_d8f4;
        state = 128'h995c_c020_9c4d_a638_ecdf_26df_48c1_f4f4;

        #200;
        key = 128'ha70c_f7a8_6f48_b367_7af3_29d4_21f4_0484;
        state = 128'he3f2_5c0f_b562_def7_6466_1fff_a3fb_c984;

        #200;
        key = 128'h46fc_169a_6174_45b1_5327_a880_0ca1_b7d5;
        state = 128'h7c83_95cc_7c94_be28_d554_781c_b691_1ae6;

        #200;
        key = 128'hdf77_fe6c_b9da_9d52_cd73_682b_6fdb_3e5c;
        state = 128'h6472_1a3f_5488_602a_2d8e_c403_4be3_851e;

        #200;
        key = 128'hda94_6f1c_c67b_3ce3_43c7_2359_70dd_350e;
        state = 128'h7c89_45a5_1e92_120f_f035_e5c4_bbc0_605a;

        #200;
        key = 128'h0084_85d8_e564_4d04_e111_11d3_8d64_a080;
        state = 128'had67_6c88_06fe_76ee_5a39_e568_84db_e27a;

        #200;
        key = 128'h174c_ddb4_1119_b017_a3fa_083f_4c07_6cc7;
        state = 128'h7172_ca39_3217_fdec_408f_bacc_e8f2_b3cf;

        #200;
        key = 128'hc57c_81d4_3871_e5e7_2ba1_0feb_bf74_df58;
        state = 128'h9d2d_05af_04a3_414a_6b00_87ff_ab8b_96cd;

        #200;
        key = 128'hf12b_b483_ff5a_cd6f_f335_f1a3_0a22_5954;
        state = 128'h775e_9b9b_f177_eff8_0b19_6003_4ac8_2778;

        #200;
        key = 128'h5886_4b8b_529a_6811_1ae7_b239_cc69_a75a;
        state = 128'hc400_5caa_2594_876d_b900_d452_6cca_a465;

        #200;
        key = 128'hb901_3da6_952f_5b9d_f7f5_7e2b_452f_4265;
        state = 128'h0965_9456_75c0_4032_5f20_fd93_c8f4_d8d1;

        #200;
        key = 128'ha5b2_1029_4bb3_fd74_28e1_6f5b_d4f4_e0cc;
        state = 128'hf184_8f05_be5c_c6d6_bb2a_2df7_32b9_f1ff;

        #200;
        key = 128'hc876_7a42_5d40_5188_52d1_b979_cf8f_497b;
        state = 128'h39bd_778d_3103_131c_6ad7_e860_89c9_1ab2;

        #200;
        key = 128'hf8bf_510c_4727_c4e0_e94f_337c_9c71_0cf6;
        state = 128'he15b_340c_3a22_086d_5ce9_e27c_bb8c_9714;

        #200;
        key = 128'hb26e_66c0_169f_e149_ce3a_1ae7_cf11_60d8;
        state = 128'h2922_4c2b_90af_c81c_0273_5ae1_d1aa_08d2;

        #200;
        key = 128'hc5e0_a7da_55af_2cd6_812e_ed79_f02a_5be8;
        state = 128'h6f5f_e0a8_2ada_5668_e4ca_0809_8474_0b0c;

        #200;
        key = 128'h5e45_2eca_e466_a024_2bd0_b9bf_98a7_d2c4;
        state = 128'h0fc9_1946_ed00_2963_207b_2777_1495_27c0;

        #200;
        key = 128'h1422_bc5e_4fa6_e7d7_0c09_4998_bbcd_adc9;
        state = 128'h3aa7_caeb_9222_65e5_b981_c385_cf2e_2620;

        #200;
        key = 128'h736f_8b59_f6c5_7d9c_5ff6_5690_9457_4d7b;
        state = 128'h7829_7d13_6dcb_b638_6beb_b62c_e79f_84f2;

        #200;
        key = 128'h08e5_6c6c_a8f6_6c63_5051_66c8_ef03_6ecd;
        state = 128'hd1e2_2c35_6c6b_87c4_6a6b_6719_236a_9b10;

        #200;
        key = 128'h5cbb_6b2f_59e4_eafc_0d08_d26f_4429_a58d;
        state = 128'h74a1_7ddf_504e_2a57_9450_1d9a_a81d_990b;

        #200;
        key = 128'h309c_948d_44a7_20d7_f05f_2f75_6b51_29dd;
        state = 128'hc84c_0b59_d4aa_ff5b_4707_179c_ddcb_4ac5;

        #200;
        key = 128'h844d_ea61_85a5_dc3f_adfd_5265_3944_8098;
        state = 128'hdd47_a513_2450_843c_1c12_8ed0_d848_f572;

        #200;
        key = 128'hcbc2_5d4d_6c1d_8b17_599c_419f_6552_7187;
        state = 128'h752e_5ea5_be3e_8a7f_3811_5b20_5b21_7f34;

        #200;
        key = 128'h4981_f34b_25ba_19d0_975d_db08_0e02_b483;
        state = 128'hbef9_61b3_a28b_4549_bf81_8f65_0534_a581;

        #200;
        key = 128'h4c09_7849_a9a4_0240_3e2f_64cf_3eea_0d94;
        state = 128'h9b0c_0a8d_8aa4_3828_e404_62a9_9cde_84b9;

        #200;
        key = 128'h1042_2df5_b69c_cb3f_e570_cc2e_3b76_cef2;
        state = 128'hb528_dcbe_b45d_761e_221d_32f8_eb04_a1bf;

        #200;
        key = 128'h73e2_b851_a39d_333a_869e_9e68_192a_9fe5;
        state = 128'hd71c_0553_41ef_4adc_79de_8279_1aa7_8aeb;

        #200;
        key = 128'h1251_a219_56e6_d998_3754_e378_b614_3b97;
        state = 128'hae09_df69_458a_3533_ad85_083f_0c77_8f97;

        #200;
        key = 128'h28ac_c9ea_696f_1ed2_3e02_7e2d_1e84_b71b;
        state = 128'hc37d_7f27_87b4_0475_2321_7e17_8593_7733;

        #200;
        key = 128'h073d_2537_c8dc_7f6a_1506_cd0a_00e6_f919;
        state = 128'h2331_38ea_4e76_74ec_4484_0b18_1dd4_c05f;

        #200;
        key = 128'h72a7_72fd_4500_a641_0800_27e2_79c6_026b;
        state = 128'h07d7_9d56_26f5_3332_27ca_0a04_f7f7_4c91;

        #200;
        key = 128'h99e8_a164_c8f8_526b_7014_b424_9fe4_0be6;
        state = 128'he8a8_bc2a_2e25_3861_dbb7_a828_6204_80ef;

        #200;
        key = 128'h5bb0_c0c9_7dd3_c636_a141_993c_34b3_1b67;
        state = 128'hd4fa_f26d_3c75_ff26_adde_85e4_b0f2_b075;

        #200;
        key = 128'h4e94_1fcb_450f_97f3_769c_dc0c_77b2_b1e7;
        state = 128'h5917_2227_578e_cbd0_6a50_5021_32c8_1868;

        #200;
        key = 128'h301b_c3d6_4a40_9058_e189_fb5a_9b85_edec;
        state = 128'h9937_11ac_a7b7_77a9_874f_6818_1537_5ad9;

        #200;
        key = 128'h198e_36f4_ba35_cefd_3444_37d6_a901_ea00;
        state = 128'h8f66_0ad8_5000_a0c8_54fb_7ee4_b108_e15d;

        #200;
        key = 128'h923b_98dd_150a_701a_7b27_c5e0_3893_7085;
        state = 128'h1caf_101a_03f3_46f0_357c_2e2d_760d_f1d4;

        #200;
        key = 128'h12ae_5ace_0f21_a0fc_481c_5267_061b_fa6b;
        state = 128'h4f3d_6a74_5e26_94eb_a710_3026_6b50_909a;

        #200;
        key = 128'h550f_9bd9_f60c_635f_2db7_d4cb_594e_2dbb;
        state = 128'h1a31_7035_554b_ad7c_be52_5a75_31c7_2813;

        #200;
        key = 128'hf3df_c0ec_5996_fbbe_8191_f0de_7e39_349f;
        state = 128'heca5_6145_b7a5_246a_5bb6_2158_db06_6cf7;

        #200;
        key = 128'h671f_2c37_01eb_b603_3bbb_fba6_d19f_2bc5;
        state = 128'hd56c_9fed_f1e3_3317_d4ba_eda0_4236_f29c;

        #200;
        key = 128'h6147_d5a5_b7ce_3fa5_a359_4a0b_af2b_f034;
        state = 128'h313f_448c_3a80_7e8c_7a5b_5dd8_1892_cfba;

        #200;
        key = 128'hf296_2760_3d39_8e77_c363_c67c_3959_3919;
        state = 128'h7139_d020_239f_cc54_19a5_764c_f45b_2c54;

        #200;
        key = 128'h0fd6_24ec_6af1_1a4f_9b36_b54a_33c0_0388;
        state = 128'h043f_1dbc_30f2_6f47_27ce_b99a_c4a0_9a95;

        #200;
        key = 128'hbef9_86bd_ccf9_32a8_fbd1_21f3_7837_9c0a;
        state = 128'h4bd1_a88c_fb2c_de32_d3cf_c88e_c13d_fcaa;

        #200;
        key = 128'h6a1d_1d27_ff2b_85d6_874c_39a7_1736_2fe4;
        state = 128'hcc38_f49b_35a6_6626_c7dd_ffd9_c26f_02a4;

        #200;
        key = 128'ha1f2_99f0_c2ce_5b42_ef90_e86f_d00b_a11e;
        state = 128'he6fc_eaa9_d520_f2af_5bf7_2e3e_ccf4_699d;

        #200;
        key = 128'h79cd_008c_9093_9c60_829a_4e2c_dfa8_c0f2;
        state = 128'hd39e_78a2_9cf7_ffb5_2829_e8a5_9204_3846;

        #200;
        key = 128'h7662_6c7a_12b6_b6b8_103a_8c7c_3e06_aaef;
        state = 128'he46c_4ec1_2c38_7639_69b3_ce19_4194_78b6;

        #200;
        key = 128'h63d3_7533_b20f_0336_61d5_6d22_37a0_6cad;
        state = 128'hf6d6_81e9_9865_e89d_93b1_b85c_f413_a0ac;

        #200;
        key = 128'h36f9_bac3_0670_ba2e_7a75_cda2_f762_17be;
        state = 128'h21a2_8b17_6d78_1ce8_a4ed_ce86_d862_4f64;

        #200;
        key = 128'h8f2c_599a_3022_964b_9957_f77c_3fc4_9e91;
        state = 128'h2aac_d3d2_f4ec_0f13_7353_49c4_d9ca_cfca;

        #200;
        key = 128'h97dc_6836_5215_422c_969e_6a36_796b_23cd;
        state = 128'h5424_4911_da97_1280_dba0_3ed3_3ae6_d7c9;

        #200;
        key = 128'h4f3f_a959_bdee_031b_c329_4e45_f4d8_173c;
        state = 128'h2b0b_7d91_c946_20b5_001c_0ad4_2ede_5035;

        #200;
        key = 128'h47ee_f857_c31f_df25_c0fc_1da8_8cda_0c9c;
        state = 128'h1580_652c_4329_3345_87f5_17f8_844c_7fd9;

        #200;
        key = 128'he4d2_c499_fe52_bb5f_0f0f_3066_222c_2409;
        state = 128'hab5a_542f_0e9b_f39a_b650_c223_bed4_c4ea;

        #200;
        key = 128'h6ba5_74ff_b25e_6fc7_3fe2_c151_1b0d_24a3;
        state = 128'h82c6_02f7_6e40_e73c_27f6_e78b_44c9_2e43;

        #200;
        key = 128'hd599_8c29_cdae_d825_1e84_c679_1b6f_4381;
        state = 128'h1e95_8c9d_6d46_7550_2857_5940_81b9_6abc;

        #200;
        key = 128'hd129_d946_322d_14ab_99cb_c1ce_20bc_f409;
        state = 128'hbb29_9d2c_15c6_ea33_3f3e_2ca9_3f05_97d7;

        #200;
        key = 128'hceec_449b_1d55_cf2e_ba9f_b92a_7896_ff9f;
        state = 128'h4a64_0da6_df1c_abf4_1154_e522_23da_ad5e;

        #200;
        key = 128'hab07_89ec_e0de_cf6c_340f_9fdb_2af7_da81;
        state = 128'h548b_e97f_612f_9745_1260_56b4_fa8f_166c;

        #200;
        key = 128'h0ab3_d9c5_8a47_7586_400e_47c2_fe86_f14b;
        state = 128'hc897_eaae_66de_8e23_bd54_2708_8885_063a;

        #200;
        key = 128'h78c2_9f90_8596_3737_812a_6343_74f1_82be;
        state = 128'h99b4_5102_784b_c51c_f3ed_1822_0eb2_7691;

        #200;
        key = 128'h4ad3_3ad0_5caf_df63_5f1c_738d_9977_385a;
        state = 128'hc967_1cfb_e9be_a580_8502_63e1_61e3_da66;

        #200;
        key = 128'h78c1_576e_a354_9437_5917_2c08_65cb_7448;
        state = 128'h7485_b7d0_36bf_f7bd_b854_0ee3_a232_6216;

        #200;
        key = 128'hca17_da07_84cb_5adf_cf74_e146_f128_7757;
        state = 128'h69f3_88f0_2d0f_5f90_fb65_b0ef_f05c_2668;

        #200;
        key = 128'h7697_12cf_79b5_cdf3_a7f3_a781_cfed_0455;
        state = 128'hf7a8_826b_896a_72f5_7e71_9b3a_e58c_5c06;

        #200;
        key = 128'had9a_5557_13b9_698f_93da_82f2_1a34_b8aa;
        state = 128'h2226_eb77_1b78_be01_00b8_0561_19c1_a660;

        #200;
        key = 128'h9cd9_754f_51e1_e366_e38f_d9cf_97db_fdd2;
        state = 128'hf570_318d_19ed_73dd_770f_c044_0594_c386;

        #200;
        key = 128'h85c0_cba1_22da_651f_7355_02e0_b28f_e785;
        state = 128'hac0a_ad82_5f57_c8fe_1c3f_6837_c8bd_b3c2;

        #200;
        key = 128'h8310_a678_219e_b741_c201_4aee_ead4_9231;
        state = 128'h9c8a_613d_602c_e0f9_f2b6_186e_8b04_12dd;

        #200;
        key = 128'h904a_77da_b0ff_1cc2_2adf_1fee_b2e5_6368;
        state = 128'ha1b2_6417_2291_6d43_4466_18fb_8964_52c6;

        #200;
        key = 128'hb01e_3e0e_8840_2ce8_6778_cec0_0148_e8be;
        state = 128'h80ba_8fc3_b24e_e196_2972_fbde_8601_7e8a;

        #200;
        key = 128'hd782_8ae1_23fe_20c4_ec2e_4eaa_cc0d_9a17;
        state = 128'h7493_0a24_58f9_ee8e_283d_9225_d5af_765d;

        #200;
        key = 128'h9c87_e45e_cabe_78ef_a529_63d2_90c4_2e2a;
        state = 128'he9a9_be3a_45dc_4c17_621c_6eba_f864_da00;

        #200;
        key = 128'hc15c_3270_ee1b_615f_a425_092b_eca8_9239;
        state = 128'h0d1d_928b_2204_db1b_e93b_7322_5cbb_3a21;

        #200;
        key = 128'h142f_164a_6f86_b366_b1a3_67e0_b9ef_34f7;
        state = 128'h7ac6_6d72_a686_b294_0f11_3219_3360_e42b;

        #200;
        key = 128'h4f0f_06ff_0bdd_fe25_4e3d_68c1_c4e2_6826;
        state = 128'h8107_58c9_7804_bc73_187e_f782_45c9_febc;

        #200;
        key = 128'hf70d_4034_b3e9_bc58_8712_7a8f_b800_18ed;
        state = 128'hb168_c7d4_655f_e4a7_f63f_fc8f_b6f0_9f3f;

        #200;
        key = 128'ha326_3feb_63e1_ceef_9464_899e_5207_0161;
        state = 128'hbe07_cdf2_2ae6_d6c4_88ef_b8c2_fcb7_92b3;

        #200;
        key = 128'h9561_f353_246e_83a4_6acb_7247_a7e1_b2f4;
        state = 128'h01a2_c468_4806_1cd6_7ce0_abb4_a94e_e103;

        #200;
        key = 128'hcb24_5d84_624b_cad9_4145_4d49_df59_d13e;
        state = 128'hfd9a_44ff_c17d_3afd_6919_76a7_3427_7769;

        #200;
        key = 128'hba72_7fb3_f494_2675_51cf_d277_af0c_0c53;
        state = 128'h34e5_e974_4b59_0494_b79c_56fd_eeeb_4bf2;

        #200;
        key = 128'hf9b1_75eb_e7b6_16f4_6fd3_b453_c465_36f6;
        state = 128'hc5ca_cafa_8d4f_bd0e_08f1_a056_6457_c87b;

        #200;
        key = 128'h4a1c_8ed9_9348_1ed6_8ea9_70e6_52b1_4ff3;
        state = 128'h1c76_2005_6438_2692_4fe9_6187_8838_ff96;

        #200;
        key = 128'h78a0_ae05_2e84_2422_d68a_b1e3_8eb3_29d8;
        state = 128'h57d3_b86e_6e1f_7b41_8b01_7c38_092b_f1c6;

        #200;
        key = 128'hc51b_0206_5b11_396f_1ee7_912c_c2dc_befb;
        state = 128'hddce_9f4d_adf6_c9fe_6083_36e3_7147_ba83;

        #200;
        key = 128'h6142_02da_b3bb_37be_5d00_8ecf_8452_319a;
        state = 128'h5a4b_8684_10fa_612f_5c3c_b185_4279_198e;

        #200;
        key = 128'h8fd0_5ab2_fa7e_fa76_f6d4_d5c4_4f1f_ae28;
        state = 128'h862c_a192_ae96_858b_82ea_8f4c_fc15_5805;

        #200;
        key = 128'h85c7_b3ff_ec61_c324_6e81_16b7_2663_4d0a;
        state = 128'hac4e_5a78_a30e_9bb8_fccc_f26f_a16f_3cbd;

        #200;
        key = 128'h11d7_5c6f_08ad_4011_c3a5_bb12_984c_56b0;
        state = 128'ha5e0_0b90_2c53_3cdf_69f1_0f0e_9b5d_41b2;

        #200;
        key = 128'h5cc3_792b_11ea_e74c_4a45_e18d_915c_4247;
        state = 128'hacd4_8f68_a2a1_0f2a_4ca0_282c_e783_5ae4;

        #200;
        key = 128'hc2b6_1e01_4aad_5398_42d4_4a8f_ee3d_f46e;
        state = 128'h06ed_1fcd_1ecd_89c6_3f8f_9865_2c1a_49dc;

        #200;
        key = 128'hee82_26df_c786_97f7_e368_e562_403a_322b;
        state = 128'hb966_4367_5b21_dfe5_7038_6654_9ff6_e797;

        #200;
        key = 128'h72fa_d787_78ed_cde8_369e_d725_b241_cdb9;
        state = 128'ha46d_2a24_6bc5_fccc_08d2_b115_abc6_f433;

        #200;
        key = 128'hc424_a794_e322_4f73_9ac9_2b28_9aff_2e0f;
        state = 128'h1ff2_e291_2f93_93a9_f3c0_83eb_6e8f_93af;

        #200;
        key = 128'h0c2e_8c4b_76bd_803d_3bcc_cad3_7d0e_e5cb;
        state = 128'h3224_f536_6b97_292c_adf3_a7cf_aed8_054e;

        #200;
        key = 128'h345d_622c_e052_6777_6fca_971e_103e_0a5e;
        state = 128'h5bb8_422d_14e5_edba_22ff_76ad_ef61_0336;

        #200;
        key = 128'hbaf3_8965_775b_0b03_b750_1aaf_9fbb_bab7;
        state = 128'hfce4_dd62_782c_8e56_28a5_05ec_02bd_30ca;

        #200;
        key = 128'h4aca_85e8_5755_c802_6899_3b60_2e8b_6121;
        state = 128'hd9fc_59cb_6012_f2f7_e41f_db33_55b5_381b;

        #200;
        key = 128'hff9c_a417_6fdb_5d38_9ed8_299b_e357_7186;
        state = 128'h2664_61de_baed_5e59_516f_c9cf_afcd_5d3c;

        #200;
        key = 128'hab58_7421_6cf6_3847_e06e_c535_9c14_84f9;
        state = 128'h3ca6_b41b_d64a_acc8_39f4_6e20_9195_4ab4;

        #200;
        key = 128'h480c_0b59_088c_5ded_ecc0_f857_6a36_6f02;
        state = 128'h9e22_621e_e705_aaed_27ed_b535_3174_404b;

        #200;
        key = 128'he3ee_d509_6601_0a70_d27f_cf48_4ed3_3cd9;
        state = 128'hd602_d0bd_8ef4_2cbb_ca00_8e7c_28fd_ebb5;

        #200;
        key = 128'h30b6_4af8_b705_4614_4e31_2470_4c64_2abc;
        state = 128'h5b6a_b019_c441_a01d_3687_b338_12b2_9b41;

        #200;
        key = 128'hc7e7_b9e7_0961_b800_5274_4d5b_1ac6_365b;
        state = 128'hb39a_2638_7711_98ba_a4f9_1b28_4f36_e2f9;

        #200;
        key = 128'h7079_9193_8ed3_0355_0dfa_a082_4c83_e0c6;
        state = 128'hec30_5eda_7474_f171_21ca_0612_8b8c_e067;

        #200;
        key = 128'h9489_11fa_2393_d31b_7553_4fd2_a8f5_f098;
        state = 128'he53f_95a3_8359_8b13_67a5_e8a0_42d3_4611;

        #200;
        key = 128'hb716_796b_2c5d_edd5_a71b_ecd8_005a_0d07;
        state = 128'h0d3e_1cd2_11fd_468b_43b2_46e8_0fd8_caba;

        #200;
        key = 128'he190_6454_46c9_0f83_02c6_c799_fa8d_fd74;
        state = 128'h2760_335f_8a2f_7dbe_fa69_1905_beec_1cc2;

        #200;
        key = 128'h989f_404a_1bcf_2472_9e2e_88cb_a326_2a9a;
        state = 128'ha0a1_0aa1_298b_e391_f14e_c4c2_a708_0c28;

        #200;
        key = 128'haa29_717f_7c57_2453_136f_b01a_d8ef_3e08;
        state = 128'h47e8_36f9_66e8_ee0b_efd7_f99e_ba50_d5d1;

        #200;
        key = 128'h99eb_6d8c_4795_ca35_099b_0a71_8e91_68e9;
        state = 128'hbe82_f815_5530_d53f_5159_6e7f_bd9b_3c17;

        #200;
        key = 128'ha809_1a64_d2d2_69e8_0ce5_96df_fc3e_f8ba;
        state = 128'h0fe8_1e12_a849_98e3_8065_8c5a_c2c6_30d5;

        #200;
        key = 128'h8d67_c892_fb99_0642_ebe1_a5f8_5b16_c560;
        state = 128'h4f2c_6de2_047d_e3a5_06bd_3a3a_3c90_a84b;

        #200;
        key = 128'h687b_6226_d09f_cf95_187f_0f21_227e_8cc4;
        state = 128'h7d45_d7ab_a612_5177_a241_4d54_ddc6_a5c1;

        #200;
        key = 128'h201d_ded1_8d5c_5981_f117_3ba1_9376_815b;
        state = 128'he53d_eeac_ca67_bce4_7912_4d37_ebe9_9e29;

        #200;
        key = 128'h6076_ae1e_f358_1a0c_210d_768e_209f_08ec;
        state = 128'h2554_eb1e_fd61_164c_e5d6_7eb7_3653_9561;

        #200;
        key = 128'h63d8_9e70_2470_03ce_8c80_6493_846c_9b1f;
        state = 128'h8608_ce0d_505f_980b_937b_1cde_0be5_3cfe;

        #200;
        key = 128'h854f_8cda_e6dd_3a71_bf08_30b0_b3bb_7a6d;
        state = 128'ha288_4cb2_811e_745b_a30c_9fb1_8da3_aaa6;

        #200;
        key = 128'h9433_5c1e_1a42_23b0_ff31_0295_a66e_f273;
        state = 128'hf97a_bd1b_b866_ed83_291e_18ad_45e8_bb61;

        #200;
        key = 128'h5604_4314_8ebe_c5df_420d_b8e2_8c57_5148;
        state = 128'he8ac_9455_6792_5ad3_8348_5602_205a_7e06;

        #200;
        key = 128'h64fc_95bf_f8b1_1444_efd7_cb04_f508_61b2;
        state = 128'h32ce_1c15_2efb_7fb9_8a54_b678_46f5_f52b;

        #200;
        key = 128'h1016_7ffb_a739_5c06_35fc_d749_ec48_6ef1;
        state = 128'h9945_91e5_e756_cb57_efdc_a744_9032_756e;

        #200;
        key = 128'h3719_6ccf_ff8f_1a66_1326_be09_0b13_3a3f;
        state = 128'hb6d6_df5f_c270_f2d5_eb43_314b_ac33_400c;

        #200;
        key = 128'hc0c1_47be_c580_5723_ac06_c1d1_05c7_1eaf;
        state = 128'h37b4_bbaa_eb91_607a_e44d_1754_5c5d_86ba;

        #200;
        key = 128'h1df6_b087_6c58_abfe_7eef_7042_c58d_8804;
        state = 128'ha8eb_bbd8_4c77_559b_9f2e_6362_7e29_7e0d;

        #200;
        key = 128'h03d9_88f5_24d1_0117_11d4_f953_0b2d_fab1;
        state = 128'he606_a424_a7c2_b1b0_1fda_d610_67d1_8ca2;

        #200;
        key = 128'h48b5_207a_2076_3ecf_239d_4060_c31d_4d75;
        state = 128'h2c13_6210_f440_6879_5af2_d88f_c9bf_0944;

        #200;
        key = 128'h66ce_37a7_e4f6_dda0_9acf_1e28_6aee_eb4f;
        state = 128'h39da_fcaa_6d35_e69a_7631_316d_b5f6_0472;

        #200;
        key = 128'h16ed_1b1e_471b_f95d_ec19_cc96_06b6_8519;
        state = 128'hcb01_c31a_9fd1_1494_98df_bda9_312e_029a;

        #200;
        key = 128'hce2b_df51_5e22_786f_bb2d_640e_0b97_0faf;
        state = 128'h7343_538d_2422_9b09_8481_e077_595d_91e4;

        #200;
        key = 128'h7353_8ef0_77e2_bbea_7b39_0d97_7724_4b57;
        state = 128'ha99e_7ee4_9435_f816_64a0_8e86_4a2b_99b8;

        #200;
        key = 128'h4174_7908_fc0c_f6d7_9b1c_b51a_6d82_a406;
        state = 128'h2eae_3833_81c7_3c90_42fe_6924_0b1e_69f9;

        #200;
        key = 128'hcaaf_7df2_4035_25bd_1d05_6470_0080_fe64;
        state = 128'ha27d_1e53_0f47_fbb8_fd1d_e65a_e66e_33c5;

        #200;
        key = 128'h057e_d5a6_e628_5feb_a35c_a571_0952_b882;
        state = 128'he310_e315_b79d_f141_d269_8315_9af8_64dd;

        #200;
        key = 128'ha762_5440_64ae_3d1e_3404_fa4a_bec3_f545;
        state = 128'hd7ca_d2bb_b45d_6261_3cb9_a08f_a255_ca05;

        #200;
        key = 128'h0e19_f40e_9f9f_a69a_c87e_b736_bea0_bcef;
        state = 128'hae64_ab4d_7636_e1ca_ad8a_d99b_12e1_1c4e;

        #200;
        key = 128'h701a_9e78_597e_5964_b96a_009c_8016_ef29;
        state = 128'h6540_6d35_0990_8ef0_0ee1_60ef_9496_7d09;

        #200;
        key = 128'h7b09_7c0d_2ae9_6461_58fb_6c8a_093a_a6a0;
        state = 128'hf2ec_7b41_b9a3_881e_ab52_2ac2_cb30_cd01;

        #200;
        key = 128'h67a0_8dc4_aa3f_7a33_c53c_769c_5e6d_ccf4;
        state = 128'hc784_b81e_f2ed_0a53_4831_3b39_fbf6_ad0c;

        #200;
        key = 128'h5bac_4466_dd10_81ed_060f_57ea_f56f_37b2;
        state = 128'hca89_916a_f5ec_0404_5187_162c_b0b5_feef;

        #200;
        key = 128'h6613_2e93_ef26_2f55_9340_9de7_1c94_e2cb;
        state = 128'h35eb_475c_ee57_b6fe_6c50_1ae1_e70a_7205;

        #200;
        key = 128'ha841_85cd_8d09_8640_f086_713c_6b49_4f3f;
        state = 128'he221_4bcb_9979_693c_63e3_0af1_5b0e_d043;

        #200;
        key = 128'h81c6_9a69_9f9a_fe3d_1d91_126e_1e2c_9818;
        state = 128'h0a95_b8ed_674f_00ea_425c_1bb8_11b4_7cab;

        #200;
        key = 128'h51d7_8750_8eda_cb80_7f39_7362_587e_fcc5;
        state = 128'hb423_cbdb_0874_ad4c_ec4d_282f_9dd0_bb01;

        #200;
        key = 128'hf090_b662_bea9_6597_9c78_f085_11ee_3901;
        state = 128'h72ec_c042_1d65_3e0f_0bec_46cd_bde7_3ab0;

        #200;
        key = 128'h53ab_9fa7_e4c8_9d81_8a85_9b36_975b_8093;
        state = 128'hcddf_cb5b_7168_9558_dec1_cda2_b250_b4bb;

        #200;
        key = 128'hd62b_013e_b696_f779_f780_4eaf_9579_4b52;
        state = 128'h1819_5541_a9f0_23dd_98c7_c54b_2fee_e80a;

        #200;
        key = 128'h682e_b75d_fa94_64de_6d99_e4a7_4e69_7bfb;
        state = 128'h7009_8087_63f3_50ca_52b2_850c_c131_9bf9;

        #200;
        key = 128'hb2af_de06_26bd_67e4_abe1_c4d8_c927_8102;
        state = 128'h5b29_db0d_0c35_c003_7bcd_5ac1_c082_fff4;

        #200;
        key = 128'h4841_c8b8_0cc1_98d1_b37e_5cd6_01ec_e6c4;
        state = 128'h17e9_2f55_5ac0_52b6_85bb_b894_d707_1e68;

        #200;
        key = 128'h49b6_50d9_7e17_671f_8b37_2300_b5ea_0ffc;
        state = 128'h045e_abb5_b123_4d7b_69a2_901e_51f0_bcaf;

        #200;
        key = 128'h17e9_f840_cb43_a568_468f_4725_3016_f086;
        state = 128'h02ec_dcbd_3a68_7ca6_0edb_d76c_9a07_9f46;

        #200;
        key = 128'h80fc_1d6b_a0ea_5da4_abad_0cf7_55f1_277a;
        state = 128'hd926_0163_ccb0_6611_a385_5ef8_dee7_0f2e;

        #200;
        key = 128'hc266_e62a_4d4c_9899_31aa_0512_d8af_3dff;
        state = 128'hcf4b_cd1a_09e1_121b_e926_3d13_eea1_224e;

        #200;
        key = 128'hb75c_24c1_224e_de8f_b81c_2ecd_912d_7140;
        state = 128'h25fa_df53_6bdc_ae4c_fef7_785b_7ff8_084e;

        #200;
        key = 128'ha167_fb5f_98fc_599b_4de2_8fc8_3f90_42e7;
        state = 128'h9101_202f_2863_0129_c068_f7de_fd46_e453;

        #200;
        key = 128'h0921_f14d_da97_c75b_132b_aa92_cc77_cab7;
        state = 128'h4fa6_bf99_0c64_f557_8f2d_708c_729a_9e3e;

        #200;
        key = 128'h23f8_e5e0_ff5e_c8e3_d595_1d85_20f0_8518;
        state = 128'h4904_6042_741b_130c_8e96_1da8_ac20_bfc2;

        #200;
        key = 128'h31ec_d709_1da9_2f25_82a5_5ea3_364e_f79b;
        state = 128'h665f_6427_af6c_19fc_a1c6_c85a_1107_f407;

        #200;
        key = 128'h70db_4333_cc3d_b2dd_6d18_fb17_b1ca_bc42;
        state = 128'h3754_3b6c_ec90_0063_61d9_3a47_1ed0_5a02;

        #200;
        key = 128'ha0cf_4ee0_1fab_11ac_d892_37f1_38dd_827b;
        state = 128'h48a6_125f_6b0c_9206_9529_3473_9474_3cdd;

        #200;
        key = 128'h2309_a953_fec8_e40c_ce81_c564_8543_6e39;
        state = 128'hd3e7_ae4b_c4e3_53bf_87e4_cca1_f8ed_deab;

        #200;
        key = 128'h024f_d907_7f61_ad9f_5166_63fb_ae3e_a3da;
        state = 128'hddc3_a7ee_d6fe_00fa_42f9_5a81_46e2_2401;

        #200;
        key = 128'h6b55_e6f1_a9eb_1ec5_d8cd_d929_54e9_7a9e;
        state = 128'hec5a_f6c1_4806_840a_6b5e_8889_ecd9_89cb;

        #200;
        key = 128'hdf1d_c5a5_f244_b158_337c_e4cc_e23f_5fae;
        state = 128'h9dea_eb45_7211_8a3c_daab_a9a0_4930_dfca;

        #200;
        key = 128'h7ae9_33d6_8ed6_f165_c083_6581_7c48_6d01;
        state = 128'h94a7_2b74_9549_04a3_d2f3_9786_58f1_9d92;

        #200;
        key = 128'h0263_0ba1_01de_9e36_e81d_9708_f3e9_8cf1;
        state = 128'hda7e_e134_bf6e_1879_f1a2_7b60_becd_0b4c;

        #200;
        key = 128'h2112_2fcf_b2bf_cab2_9912_d8f9_7f49_39ac;
        state = 128'h263a_96b9_5243_9096_6d78_59ef_d1f0_db7f;

        #200;
        key = 128'h0056_8522_2ac1_d0b3_4ae8_6ded_9e8b_eff9;
        state = 128'h091b_299f_3129_4054_cf4a_c46b_abfb_16b3;

        #200;
        key = 128'h9c94_a6b1_ae65_335a_0a52_d42b_7d1e_6062;
        state = 128'h57d2_3e21_190c_7453_cbf9_57c0_7cb2_1ed9;

        #200;
        key = 128'h9610_1d0b_2b66_7a9a_5477_a417_4abf_b30f;
        state = 128'h85d1_96c4_9cae_00ca_4a87_872b_edcc_f010;

        #200;
        key = 128'h6b4b_34f0_3190_80fe_c6d8_2ac4_b8f6_70d1;
        state = 128'h0815_932e_c961_2e33_6afd_272d_970a_3b43;

        #200;
        key = 128'he370_2d63_6228_e5e3_7b10_66fe_1f46_70b9;
        state = 128'h7045_8808_82c6_552d_0e15_b936_5bf7_294b;

        #200;
        key = 128'h7851_87e9_3663_8709_e300_d5f0_169e_33e5;
        state = 128'h2a58_7620_e58a_0041_5330_e3d5_caa1_d1f6;

        #200;
        key = 128'h3490_958c_9081_59e3_9387_75ab_e3bd_2f85;
        state = 128'hb997_cb99_e850_21ea_34b3_06fe_5482_e9e0;

        #200;
        key = 128'h727d_d505_1b24_8d5b_b2a3_0909_7cbb_6851;
        state = 128'h3be7_78be_bc88_e7b0_66e8_ef62_3ca9_ce40;

        #200;
        key = 128'hc4fe_cff8_ccf8_babf_1ceb_10d3_4f89_4515;
        state = 128'h9447_f35c_792f_7cfb_0eab_f578_7d2d_310b;

        #200;
        key = 128'h5e74_8e74_1544_ad7a_bf5f_4602_5899_7fdd;
        state = 128'h88da_074b_f22b_1fea_16c7_901e_fb2b_e9c6;

        #200;
        key = 128'h258e_2e4e_ee3a_c965_5d67_8cbf_0ab3_6acb;
        state = 128'ha3ac_1fbb_37bc_14f6_18bb_2b02_8d5b_a7dc;

        #200;
        key = 128'h5843_e416_bc82_ac4a_0dc9_4196_ed4f_2c48;
        state = 128'h63b5_62ef_1407_d322_afe1_8e77_2115_dc46;

        #200;
        key = 128'h763c_88d7_f979_c963_c5c2_1846_a690_c185;
        state = 128'hc702_799d_13c4_55ad_016a_d5f6_3331_cf58;

        #200;
        key = 128'hd3f3_99b9_5474_b739_4a50_ead8_5774_5f98;
        state = 128'h258c_b74d_2780_9e0c_179b_5bb7_1f3d_61ef;

        #200;
        key = 128'hcf06_92c8_3c32_f20c_a1a2_4913_3046_b671;
        state = 128'h51da_dd09_b55f_07a4_a86c_b3b1_f819_5b00;

        #200;
        key = 128'h9ab3_16ca_476b_0827_3a77_a20a_a382_bca0;
        state = 128'h6b02_eb87_0f1d_21e9_e7c8_56b5_f98f_90dc;

        #200;
        key = 128'h4fc7_2ae1_90d3_bf41_b0cb_9ad4_e1e8_2d54;
        state = 128'h9d0f_29c7_58d1_74ad_5964_cf9a_360f_d75d;

        #200;
        key = 128'h8485_1773_2eef_7cbe_3deb_bd21_146d_9945;
        state = 128'ha406_1674_7dd5_5926_1b01_3320_f6f6_4523;

        #200;
        key = 128'hc582_4538_5557_a42e_e79f_7f3a_851c_5cf6;
        state = 128'h4f26_dd0f_325a_8154_81f0_3879_f69f_a51e;

        #200;
        key = 128'h84e2_c5c3_c4b3_8af9_b1b8_bec3_35d2_4eee;
        state = 128'h9276_e810_bdee_6a12_aa6f_9191_7d2e_09dd;

        #200;
        key = 128'hf0de_503f_3b99_523d_378e_85b1_3fbb_4451;
        state = 128'h1aa5_5f9e_1b86_4fe1_5e0b_70cf_9f40_be22;

        #200;
        key = 128'h6703_63fd_27a8_ba14_75a8_1c11_8886_096e;
        state = 128'h83d8_a29d_d81d_f5e9_3069_3462_bf76_c5a6;

        #200;
        key = 128'hea38_ef41_f827_6ac8_7842_d096_859b_63c0;
        state = 128'h91b7_92c0_c73e_5f3f_6d57_7e2f_e43a_f3f7;

        #200;
        key = 128'hc8cd_4366_f2d3_7440_454f_af61_2da2_8c4b;
        state = 128'hf7eb_482f_6af8_39e5_5843_f83b_a5b9_5e03;

        #200;
        key = 128'hb3ff_c1ec_9488_a524_405b_3de4_508c_9516;
        state = 128'h34bd_fad9_17f2_0011_92f5_b38d_4b7d_e47d;

        #200;
        key = 128'h268e_0785_0f07_75b5_be7b_5d22_640d_165f;
        state = 128'hb04f_276f_8810_ecaf_0c89_ed57_d600_777d;

        #200;
        key = 128'h20d9_32ab_b4fa_ff46_f397_425b_7faf_f159;
        state = 128'hde94_9d24_e0e3_5b10_bd2a_b37f_d390_f0bf;

        #200;
        key = 128'hc46d_3ba7_9f26_0900_355e_7d59_0b69_5612;
        state = 128'h3146_055c_0815_f5a5_7b59_46f9_a315_d2d3;

        #200;
        key = 128'he8e6_3fca_01ea_167b_c60b_4c31_730b_8f0e;
        state = 128'h86bd_7008_5373_6124_df12_2222_7dec_1b6f;

        #200;
        key = 128'hb7ff_abc6_d155_d117_4220_e213_0ad8_15d2;
        state = 128'hfaf4_d842_f9b5_a15a_5195_e2ec_bbb4_cb2a;

        #200;
        key = 128'h3dc5_0e8a_e0e3_8078_86e2_4db5_e6f9_0e69;
        state = 128'h0923_7db7_464a_b4cf_543a_1da1_46d0_f1b7;

        #200;
        key = 128'hcdaf_00ff_62e8_167c_87cf_7cf7_7b8b_d933;
        state = 128'h375f_8b45_f351_6d6f_a470_ab16_628c_0e3e;

        #200;
        key = 128'ha1ef_f394_bb34_c909_e631_08ab_0c26_56de;
        state = 128'h339b_506d_6f9c_d493_18c7_80b0_a48f_377e;

        #200;
        key = 128'hb025_e85d_3d27_728c_b64f_b237_770f_25ad;
        state = 128'hb8ff_0230_4ec9_f34d_ca4f_5b88_4df5_6a0c;

        #200;
        key = 128'hcede_c7cc_ead8_ff62_4634_8b49_99ad_6468;
        state = 128'h6029_306e_7c95_8198_ae28_ca09_2de2_1eb9;

        #200;
        key = 128'hebd2_23cf_7ed8_d1d3_cba0_a090_b2cd_fffc;
        state = 128'h4e69_c0f9_5e45_042f_5b2c_9f38_7e2a_47bd;

        #200;
        key = 128'h1db8_aa79_f91c_1a1f_f077_eb73_b373_a8b0;
        state = 128'h1123_167d_6a1f_d462_8168_3500_c98c_87a3;

        #200;
        key = 128'h6907_7948_664f_0f0b_7a18_9296_1d79_c330;
        state = 128'h0e44_9b06_c9fc_8dfc_161e_9eec_2141_5816;

        #200;
        key = 128'h718b_10fc_c163_d780_9947_fda0_139f_5697;
        state = 128'h76d4_645b_7628_1353_0648_cc3c_4ab3_d9b0;

        #200;
        key = 128'h851e_ddf2_38d3_cd6c_e31f_ab5b_1f45_3520;
        state = 128'h2e63_71ac_52bf_fc8b_637a_ed18_0d5e_c48b;

        #200;
        key = 128'he3d8_7591_4811_6e07_c31a_d86e_efee_8ae9;
        state = 128'hb341_5c8f_2e88_0c13_62e9_9dcc_c253_3470;

        #200;
        key = 128'h90d4_7aa2_ba27_105f_e93d_bbab_3854_e34f;
        state = 128'h694e_6111_7ea8_76ae_ee46_58eb_b4a1_86ec;

        #200;
        key = 128'h3d93_b83e_2cda_27c8_3f5a_79b6_f81a_e5d5;
        state = 128'h8eec_a581_ef21_c8bf_90c9_abb2_def5_9988;

        #200;
        key = 128'h18b9_7776_89ad_1ae4_023a_c82c_f197_cdd7;
        state = 128'hb150_92dd_bace_41c9_6d1f_a505_91df_a4ce;

        #200;
        key = 128'h2ecc_b699_f5a5_af06_327b_4b99_f879_3029;
        state = 128'h5745_38dc_481d_6c5b_1fe4_5b11_9d0d_710e;

        #200;
        key = 128'h8d7f_3c8f_4a80_d3fa_3616_16f7_70ad_c0f1;
        state = 128'h6001_aaed_30c9_0eca_4ed0_b739_6d01_ad01;

        #200;
        key = 128'h4639_4463_f219_771b_54ba_dbdb_4ef0_7b6b;
        state = 128'h2c32_d10f_e901_4093_cbf2_d7e1_b982_874e;

        #200;
        key = 128'h496b_d3c4_9722_a9f9_eeb7_82bc_f622_5965;
        state = 128'h847f_f21f_79ed_c5fa_3622_38d6_3a81_9ee9;

        #200;
        key = 128'h36e5_dc60_efaf_b041_807c_d03a_fad9_e044;
        state = 128'hd18f_c784_ee8a_1507_d41a_ff8b_1647_5039;

        #200;
        key = 128'h946f_800b_d178_6bca_eafb_3e7b_443c_c613;
        state = 128'h4d16_0687_771f_8d6d_b96c_b9e4_b378_bbbf;

        #200;
        key = 128'hbe27_acc3_b35b_b9ba_26db_29bd_4189_f6c4;
        state = 128'hdd42_8df3_10f9_4497_4a87_a3e3_e145_f338;

        #200;
        key = 128'h2c0d_fd32_d5e0_fda5_1e07_a56d_720b_6e00;
        state = 128'h87ad_6429_206c_9df1_2f8f_095f_d967_d280;

        #200;
        key = 128'h4ded_d0c4_e78a_d473_639a_54bb_b055_11e7;
        state = 128'h1ab4_aab3_89e1_7c66_8cc6_9a89_3049_9739;

        #200;
        key = 128'hd73c_8daf_fec6_0a59_a1bc_3fa2_10ec_f19e;
        state = 128'h4c42_0007_8cc2_7ec6_ec96_79a3_6c9b_6ed0;

        #200;
        key = 128'hde50_3b38_3d9f_5b06_b10a_39af_83b1_190a;
        state = 128'h67e9_dd92_cd07_af24_7c97_4f2f_98c3_d9aa;

        #200;
        key = 128'h6091_fd9d_7e95_46a7_d4b0_c485_b57c_d91a;
        state = 128'h39e8_1448_0511_ecda_2d96_d84b_c523_aabc;

        #200;
        key = 128'he809_bf2b_efaa_0e63_19a0_b92c_9c8f_1cef;
        state = 128'hf7dc_8b15_e336_249e_2d92_6b22_fa2c_b3df;

        #200;
        key = 128'hcf57_72c0_a260_3841_9024_eb8b_b24a_4ae4;
        state = 128'hc85d_a309_03b1_d3e6_e03d_20db_4e9c_f007;

        #200;
        key = 128'h1e52_49ba_04f1_3cc3_c051_a4d0_7203_c1c7;
        state = 128'h2701_11cc_ee35_0e72_7e78_ddc1_6910_c856;

        #200;
        key = 128'h89c3_a1c3_a398_3ab3_c8a2_afbc_a00c_d0c2;
        state = 128'h49b6_e01a_b14d_fd09_273e_d95f_a532_002b;

        #200;
        key = 128'h781a_18b8_7d88_137a_5857_8d39_a9f9_397e;
        state = 128'hdf6d_b980_6b8e_ff24_3c3e_8908_8fff_0c37;

        #200;
        key = 128'h1a64_3206_7ac1_d83e_938e_4369_3f6a_00a5;
        state = 128'h2dca_66f4_8487_42b3_61b8_70a6_572c_d7b5;

        #200;
        key = 128'hb466_d945_4b76_a834_cd16_1b0f_bf89_2a19;
        state = 128'h5743_3443_5bce_a8d7_f41c_774f_85b9_5550;

        #200;
        key = 128'h0704_6318_3308_ec8c_9c84_bc06_c42e_58c5;
        state = 128'h34eb_dbc0_d0ab_128a_ed7e_65ae_8a23_7579;

        #200;
        key = 128'h304f_4e65_c8a1_964f_2ef7_3c51_66c5_4e1c;
        state = 128'hf413_b5a6_8c6e_7c79_c233_08fd_5855_aef8;

        #200;
        key = 128'hb812_2e70_1890_c2f1_4c63_59f3_5045_d6ab;
        state = 128'h8c71_6629_b03c_0ca9_f30b_b272_e714_a842;

        #200;
        key = 128'h866c_db99_1927_8829_f564_d1cc_8b76_d172;
        state = 128'h86e8_313c_8631_79f5_50c8_f2c0_5830_7bb0;

        #200;
        key = 128'hd0de_412c_a55e_c42e_7b81_fc88_a314_d1cb;
        state = 128'h58e2_f8bd_5472_f5e4_4f71_518e_80f3_ea48;

        #200;
        key = 128'h4039_737b_e7e2_93db_f55c_d489_116e_1e5e;
        state = 128'he791_d333_d69c_9d29_e4c7_9871_f921_6232;

        #200;
        key = 128'h780e_dbbe_e40e_8017_428c_a831_7a00_4abe;
        state = 128'h6afc_b522_0a7e_3cab_7bbb_fb2e_6aa5_c778;

        #200;
        key = 128'hc2df_5a73_b618_adb5_4ad9_98fe_e712_9cf6;
        state = 128'hb52b_5bb8_a189_b276_bc52_679c_937d_7a39;

        #200;
        key = 128'h2eb5_6346_78c7_2414_c302_b2d1_47e5_ea29;
        state = 128'he91e_991e_1527_d00b_b8dd_773e_5199_220e;

        #200;
        key = 128'h58bb_7db8_0bcd_609e_e511_fa1b_f91c_b829;
        state = 128'hab9c_9cb8_cfa5_eb91_5ec9_3049_c9be_6982;

        #200;
        key = 128'h9af6_70c3_9460_8dd8_9579_8ea6_4103_5ccb;
        state = 128'h89e6_63c5_3290_4373_103c_09ae_3a4a_0a70;

        #200;
        key = 128'hde10_7687_7193_8d05_8e93_a772_2589_8ba1;
        state = 128'hd174_9bd2_514b_fe44_3ad3_2786_d0f8_59ab;

        #200;
        key = 128'hbd3c_6623_0dc0_dff5_1936_91ba_9300_c066;
        state = 128'h709b_e822_55d9_145f_c4ff_ff32_f8d3_2c2c;

        #200;
        key = 128'h094d_6cc6_e497_6333_a6d3_7177_6aa4_1a6e;
        state = 128'h2acb_5063_505f_f56c_e69c_3837_ef74_f426;

        #200;
        key = 128'h777a_fbc6_0eb9_1bf7_7c6c_993c_72ec_6283;
        state = 128'hc507_90af_b2a9_2b72_7a55_0962_289a_2c19;

        #200;
        key = 128'h7440_f829_f447_19a1_52f3_7ae6_4f6f_29c6;
        state = 128'h3253_1cdc_aebc_0df4_9514_1228_1b89_4004;

        #200;
        key = 128'ha092_0b9a_8274_2468_b664_f17f_f893_281a;
        state = 128'hc0c9_6b54_569e_7646_96fe_d699_d45f_fe01;

        #200;
        key = 128'h2e9f_b7c9_5146_5cf3_9a60_acff_0f33_9483;
        state = 128'h48e2_7705_7f4f_9f7c_6233_09db_5bf7_f3c6;

        #200;
        key = 128'h8a2b_7590_44a7_e5ad_149d_eb37_9c0b_c420;
        state = 128'ha72e_6869_e215_ee76_f3a4_c78b_f6f8_96fd;

        #200;
        key = 128'h488a_415e_8465_e339_01e3_3511_e125_4d45;
        state = 128'h8b06_b8e7_3196_6e3b_4ff2_899a_8612_e646;

        #200;
        key = 128'ha05b_7929_08eb_8955_bb2d_4384_ebb0_0737;
        state = 128'h7727_be4d_6c2a_e18c_fa1d_8037_1c52_8445;

        #200;
        key = 128'ha6b6_d0b4_fb06_45d8_657a_a38f_01d4_f675;
        state = 128'h0551_3243_e5d5_d3bf_0653_03ee_3f98_c103;

        #200;
        key = 128'h00cb_8336_9037_4b90_e267_6756_bfe0_766d;
        state = 128'hb3a5_9bef_3ae7_0101_438e_815d_f3e0_eef8;

        #200;
        key = 128'hbbf9_3d96_f61b_b24d_3ba4_25ce_eb89_e7f0;
        state = 128'hf413_5566_aad8_4612_4b4c_d647_4235_ce15;

        #200;
        key = 128'h29f2_e9ba_9f36_8a5f_bc34_1543_f610_2739;
        state = 128'h4ad1_2e8c_6169_0670_578f_2673_e9fa_34bb;

        #200;
        key = 128'h03b2_e12a_79ea_9da7_1c19_9897_aab0_e012;
        state = 128'h1c87_9f08_5da5_6f00_4a70_029b_c61b_26ad;

        #200;
        key = 128'h35eb_7f9c_bb47_12a6_a751_e6f0_8f6e_9daa;
        state = 128'h3da9_5114_6299_42e8_ef48_ffa8_9769_e3a6;

        #200;
        key = 128'hbfcf_0eed_45ef_50f1_e9a2_477c_f24a_c389;
        state = 128'h0916_8300_c8c4_e1f8_4999_e3a3_0939_bfcd;

        #200;
        key = 128'h5dc5_2039_3448_f70f_dcbc_9e36_fd59_a5e5;
        state = 128'hf418_19cc_565d_d7eb_0c17_09ec_056e_bc01;

        #200;
        key = 128'he352_5cd1_9dd5_f43c_8ba4_b568_b98d_1bfa;
        state = 128'h944a_292d_b4c0_ae5d_2662_4de8_e078_e815;

        #200;
        key = 128'h64a8_fc11_a38e_624a_ab8a_ebf8_690d_58e4;
        state = 128'h7dcb_9185_9e87_b79e_3408_1f28_2064_f10f;

        #200;
        key = 128'hfbc0_4c29_6e17_fbad_b80f_bb35_388a_2b93;
        state = 128'h39a9_25aa_52cf_fc91_17d8_bdc4_cf57_9d1c;

        #200;
        key = 128'h5991_3c07_11a0_257f_1a9d_c0a1_74bf_4e4f;
        state = 128'h48d0_140c_ec9e_733c_fb3f_9484_7ab5_9173;

        #200;
        key = 128'h1dd4_1932_a796_295e_1eab_4619_d4a2_34a1;
        state = 128'h9c2b_49fc_b779_6e35_6b94_ef3c_570c_7abf;

        #200;
        key = 128'h547f_845d_48fb_79e4_feb6_ed78_f0e2_7768;
        state = 128'h4417_52c9_4d8f_efa4_01ab_9861_7591_ff49;

        #200;
        key = 128'hfaf6_6428_6ba0_f5d7_1f28_8fd9_d6d1_d41d;
        state = 128'hcebb_80e0_6250_04cf_e197_96ae_baa2_61ff;

        #200;
        key = 128'h9795_14c9_41ee_3f71_2c79_1f6d_fb10_7b50;
        state = 128'h3524_c4b9_5d62_8659_2878_0b26_798c_d6c7;

        #200;
        key = 128'hfc89_859c_6646_9949_eaec_85c6_ebfe_6a81;
        state = 128'h9a17_8163_4db1_349e_4c13_7164_9dc9_647b;

        #200;
        key = 128'h768e_bb31_2ff5_03a6_c0f9_1cfc_fb59_39e4;
        state = 128'h3c0f_682b_fe93_8198_e0ae_87d7_f1c9_7d6e;

        #200;
        key = 128'h95d1_38ff_d7f9_5fcb_0dc6_fc86_8f09_a2b5;
        state = 128'h5c6c_77b5_1887_77a0_0390_e908_9f4f_f7c1;

        #200;
        key = 128'h01ec_efcc_ac08_ea46_3ffe_b342_f65b_1f42;
        state = 128'hc592_0090_972e_3e2f_c72a_6552_a7ae_beb1;

        #200;
        key = 128'h8300_73e7_f124_f125_eb59_c0c8_8acd_a626;
        state = 128'h6954_56b2_3acb_2555_bc1d_a51e_4a04_bd3d;

        #200;
        key = 128'hc1a6_d677_28da_893f_36fc_edd3_3a84_9fdc;
        state = 128'ha7f3_724f_9eb0_131d_5b03_7018_9823_a59c;

        #200;
        key = 128'h9ad8_cb07_e827_657c_fc3d_7ed2_37a6_8087;
        state = 128'h001e_8b78_44ae_7385_361f_94be_1a6f_6d55;

        #200;
        key = 128'h31a0_f076_030e_799a_5265_8264_c2f7_6e98;
        state = 128'hd291_af22_708c_2e28_8032_7613_15a6_fcc5;

        #200;
        key = 128'h65d3_51af_f1be_e4df_4620_997e_d2d4_79d0;
        state = 128'hb79b_9f9d_ca76_e2de_4954_ebf6_032f_ae78;

        #200;
        key = 128'h9e94_b7ad_acae_0d4d_5456_9db0_ac82_d8f8;
        state = 128'h5194_7ccf_c003_e7dc_7d71_e535_178c_c6bb;

        #200;
        key = 128'h00ed_6e63_224e_d615_bfcc_3ac9_989d_5d67;
        state = 128'h6b26_27fb_2d69_5d21_7fb7_09ae_7683_0365;

        #200;
        key = 128'h21a0_684d_629c_2b79_66df_1813_aae8_de1e;
        state = 128'hc0bd_720a_63cc_92d9_38b1_c4d2_bd9e_553a;

        #200;
        key = 128'h2756_9c38_dce0_644f_775f_0e52_0a36_cad1;
        state = 128'h8093_b565_24f6_5e23_0db4_4190_77f2_8eb9;

        #200;
        key = 128'hfb2d_39c2_feca_ce25_68f3_136c_241e_27e8;
        state = 128'h0da0_33b0_67bb_c195_e688_b04c_205d_1c8b;

        #200;
        key = 128'h8715_8790_593f_1918_ddeb_01aa_8f25_ce61;
        state = 128'h38b7_9a23_7449_7036_2bab_d358_354f_610c;

        #200;
        key = 128'h5e6e_8099_6ff7_e77f_3a17_5045_14ae_d3c9;
        state = 128'h5154_19e9_52e8_47d9_8621_5f90_5a83_bbf0;

        #200;
        key = 128'hc294_f634_c913_9ba1_5ef4_efcd_916c_a82d;
        state = 128'h76d4_d48f_c56a_cbb4_7da7_ec02_4627_9809;

        #200;
        key = 128'hc00b_aaf1_9dfa_9daf_09e1_cc4b_e421_e73e;
        state = 128'h2015_4950_a9e6_231b_31d5_e45d_fe68_043f;

        #200;
        key = 128'hac37_ea58_52fe_010b_af17_4ccd_c948_6a09;
        state = 128'h8e42_c860_bf44_a58e_d4f6_fc2c_c9da_f0b1;

        #200;
        key = 128'h6205_58ce_565c_fddc_7e62_aa45_0b99_9958;
        state = 128'h59a1_4bfd_21c9_bc9f_84ef_d949_2294_4a51;

        #200;
        key = 128'h6ec1_9308_d09c_3418_d16a_55bc_0bc9_9703;
        state = 128'h5a3b_a603_0999_f234_0646_2e4f_e2de_062b;

        #200;
        key = 128'hc088_3fb5_81ba_7f8d_f93f_81a1_bc0e_d264;
        state = 128'hd4b8_3fb0_42b4_82fa_c00a_29ac_c2d4_7391;

        #200;
        key = 128'h1660_c304_86a8_5904_03e0_0f38_d9d9_afc1;
        state = 128'hb292_272e_2fd2_3490_065e_4764_f8cf_f7d3;

        #200;
        key = 128'hee3e_5be0_29c9_b949_2b89_aec8_0d3b_7053;
        state = 128'h7f5b_87fe_b3f4_2a3f_94b9_f625_5397_cf69;

        #200;
        key = 128'h95bf_f476_9635_ee71_cfbf_750f_8ed5_a8dd;
        state = 128'h8d8e_c34b_39b7_8b29_5883_9449_d998_f0d0;

        #200;
        key = 128'h1a9a_451d_b054_074c_2eba_414f_fd4b_a9e4;
        state = 128'h16d2_dc67_23e8_29d7_f7fc_1bd5_4ab7_2555;

        #200;
        key = 128'h59e7_e6b6_7656_e2ca_dad3_91a9_b260_1d6e;
        state = 128'h8634_4eab_6eb3_82db_9d9d_bd5d_c42c_e4c5;

        #200;
        key = 128'hea18_4941_5883_b1a2_26c2_3ab8_c043_5202;
        state = 128'h3976_0b57_9683_fd5b_a9de_fd34_2871_b6fe;

        #200;
        key = 128'h4791_25f4_66ae_3bb8_e969_964a_74d2_cda1;
        state = 128'hb469_5bdd_e088_cd6e_771b_00de_976e_182c;

        #200;
        key = 128'h9045_ffc1_fc70_5b89_33ca_c08f_0c4c_3344;
        state = 128'h1577_1c20_383f_0707_f140_37dc_bdbf_48d4;

        #200;
        key = 128'h48ef_25a8_cb7f_b610_a05b_aa08_eed8_e499;
        state = 128'hae54_a94a_4350_3e93_444b_ee0e_ddec_dd8c;

        #200;
        key = 128'h29e7_bab1_223c_8fb5_ff73_ff6a_4d99_f8e2;
        state = 128'h1fdb_97c8_ffcd_523b_6bc3_557c_7fca_c9ee;

        #200;
        key = 128'hdc15_da35_0448_9f11_8c99_ce57_de82_7d6a;
        state = 128'hefbf_6727_97f1_18fd_0d66_c990_3b6f_5ce8;

        #200;
        key = 128'hef2a_3a8d_91e3_1622_b6d2_185d_296b_0804;
        state = 128'h096c_8279_b908_82e8_d205_00be_fa95_a68e;

        #200;
        key = 128'h6e66_5d9a_35e0_bdae_1cda_f5a4_84c7_1940;
        state = 128'hebbd_fb88_105d_e70c_d5cf_9118_6862_5ec2;

        #200;
        key = 128'hb71c_c690_a121_76c7_8d41_d087_84b9_8d58;
        state = 128'hb746_3189_eb54_c1a7_a49b_3a5d_8a2e_f332;

        #200;
        key = 128'hfd54_1afb_69ea_5638_0836_76ae_af25_e53b;
        state = 128'hebe1_0283_ca43_3e6d_6d5c_9e93_e611_1076;

        #200;
        key = 128'ha695_092a_7a7f_0098_34b9_c531_bcb7_dcb1;
        state = 128'h6531_1595_1732_1f58_d614_87ab_2a27_8ee8;

        #200;
        key = 128'h5e97_c43e_298e_6f0c_74b5_acfe_5a61_163d;
        state = 128'h640b_09c6_2cb9_964f_14e4_2497_05d9_943c;

        #200;
        key = 128'h4bdf_9c47_28d9_f749_eb38_df3f_d10e_7692;
        state = 128'h979b_84b3_cb62_ce75_a615_315c_daf9_a03a;

        #200;
        key = 128'he684_c91e_9626_a01f_bf87_0fbe_49f4_ddf7;
        state = 128'h66de_dc9b_f761_3b56_44ad_8478_c912_6c06;

        #200;
        key = 128'hd91d_6a2a_0ddf_44e4_8c96_8cbb_e4cb_2555;
        state = 128'h2f09_56ac_a1b4_ef0b_5d48_34f3_4799_7e18;

        #200;
        key = 128'h6712_ad60_3b6d_a643_dfef_8a07_1a8f_4f30;
        state = 128'h5ded_b404_1195_52aa_b6e8_0374_01b6_af1b;

        #200;
        key = 128'h81c3_0068_13f5_1797_4caf_8a7e_2181_2826;
        state = 128'hdcb9_55d3_63e9_be49_ba94_69e8_95e3_208f;

        #200;
        key = 128'hc73f_b29a_6200_f1e9_8b60_ede1_887f_d0e2;
        state = 128'hc7ea_33eb_71a6_4819_3420_a05b_e8d6_aa5f;

        #200;
        key = 128'hb5f9_2c12_5669_7c66_ed05_e043_d80c_f430;
        state = 128'h88df_4e24_0307_247c_0b08_87c8_330f_9c4e;

        #200;
        key = 128'h9143_bb99_a9f4_4f64_ed88_8705_11b6_0bfd;
        state = 128'h4fac_56e8_97dc_3aab_0ed9_976e_cfbe_5e9d;

        #200;
        key = 128'h2257_aa7c_5cab_5fdf_be97_ca40_f182_e17a;
        state = 128'h8023_d2ed_3ef5_738d_e8f5_31e5_272b_6806;

        #200;
        key = 128'h18c3_8935_8c4b_fcc5_af7a_bccd_74f6_c089;
        state = 128'he3fc_a2fa_31a9_1ce4_6c24_6b51_d65e_a8a1;

        #200;
        key = 128'h2076_da22_3547_d5bf_695e_d74b_49c4_8c3d;
        state = 128'h0c4c_47c2_97d9_64b0_f4c0_0435_6da7_1b06;

        #200;
        key = 128'h36d6_a85a_a64e_1f4d_91d9_1fe5_48a2_bbd0;
        state = 128'h8247_1b8d_93bc_efe9_11de_c244_b66c_6ff7;

        #200;
        key = 128'h9d3d_c35b_b00c_86c2_fa1a_3527_b222_3ca4;
        state = 128'hf854_3eb9_58c5_15da_8625_5952_8865_a746;

        #200;
        key = 128'h97ce_c669_f8a5_ac00_55a0_801b_5d3d_6d41;
        state = 128'h90a7_904f_6184_c4c9_85c2_244a_8351_fbff;

        #200;
        key = 128'h3d03_a4b9_d444_9e8f_73c2_2263_cd60_7412;
        state = 128'hc4ce_3d2a_8111_8a08_5c4f_ea8c_5a8d_e32c;

        #200;
        key = 128'h082a_9810_1a4e_b30a_a98e_6fb0_f424_2dde;
        state = 128'h3449_6d03_f8fc_c628_4e66_b0f2_20b7_738b;

        #200;
        key = 128'hef4f_4eb8_03df_3500_3ffa_9782_8f77_efee;
        state = 128'he400_071e_0121_6787_d324_0a4f_9b01_1406;

        #200;
        key = 128'hf7a4_bbe7_f5d7_8f08_7843_f0e7_9751_6710;
        state = 128'h7fb8_a004_444e_1e56_e2ce_d7f0_34dd_8e38;

        #200;
        key = 128'h2618_527f_ea78_c9be_bf1f_03c8_30a5_7401;
        state = 128'hf80a_8c0e_2652_c5a9_0620_31f6_37de_5766;

        #200;
        key = 128'ha708_13b4_a980_0946_9864_d35b_c71f_c30c;
        state = 128'hf3bc_bb7c_8ecf_16fd_1175_32f4_b68c_0684;

        #200;
        key = 128'h92e3_759c_1f40_6b35_cd74_d532_5125_2940;
        state = 128'h3c94_f4df_dee6_89ee_8576_867f_6129_cf0d;

        #200;
        key = 128'h9f2d_d4be_cb66_ebec_742c_11e0_5edb_b5f7;
        state = 128'hff71_6de2_3d7e_6948_d2c8_8db5_10ef_3c0e;

        #200;
        key = 128'he377_712f_aaa2_596b_3545_bec1_cec0_59b4;
        state = 128'h8158_79c6_f0d1_ca55_151d_ebd3_5e94_3c54;

        #200;
        key = 128'h1ece_2d20_938b_76cc_4f5d_b404_995a_45fe;
        state = 128'h5f53_e923_a0d6_02d3_91e6_5dde_83a7_862c;

        #200;
        key = 128'h92d6_878c_913b_d142_2fe9_d7ac_b964_c1d1;
        state = 128'hfe13_f74e_2e62_aa4e_efb3_225d_e267_f2a7;

        #200;
        key = 128'he6a4_6ed6_c9e7_2758_b757_94e5_a7ab_1552;
        state = 128'h95f3_9395_733e_2d8b_d8e8_018f_d6e0_dc50;

        #200;
        key = 128'h6836_a5b9_01be_2b08_f532_0664_3310_aa7b;
        state = 128'h371b_5dec_9110_d71a_3837_41e2_f9cb_27c3;

        #200;
        key = 128'h17a7_85a2_6c65_c560_bf8b_6aef_0caf_7beb;
        state = 128'h845c_77f6_f6e6_6f04_c068_3f60_abd6_a5ea;

        #200;
        key = 128'hc21e_99b8_3058_b475_5e9d_1320_175d_5fa2;
        state = 128'h931a_65e8_76f1_5392_7ce6_ee6c_86ef_7ab6;

        #200;
        key = 128'he105_1e13_f64b_a2d7_fca9_6f30_5c43_5997;
        state = 128'h437b_f763_5549_37f0_19bb_3f6e_ea21_a23f;

        #200;
        key = 128'h9ecb_5e3d_5335_1644_892a_9dd8_8274_349c;
        state = 128'h776e_e53c_0627_1f42_37ca_07d7_a279_40dc;

        #200;
        key = 128'h3fd6_1783_da95_22e9_f622_82b3_fa20_8bbd;
        state = 128'hfc82_97d9_36be_2d7a_f0c9_4174_0efe_6f52;

        #200;
        key = 128'hd358_c91e_387d_15d9_abee_09ee_04d8_05e9;
        state = 128'hd2d6_90f2_b500_5783_61c7_5b1d_92c4_1ce0;

        #200;
        key = 128'he016_47b7_2c33_6887_25d4_7402_c70a_915a;
        state = 128'h1d06_324e_3ebd_bad5_9a6b_2ded_23b7_d488;

        #200;
        key = 128'h6f29_87f7_cdbd_46a8_3582_324a_eadb_e3ca;
        state = 128'hc4d2_fd9b_b3f0_1600_c297_0354_68e3_b52d;

        #200;
        key = 128'h2fe6_d9cf_c190_14c0_e5e4_7338_8fba_9c26;
        state = 128'h4d73_ef6d_380e_17c0_f609_e802_14de_ab2e;

        #200;
        key = 128'h1760_5b91_9872_65fa_f9d4_1fc8_bec0_5ade;
        state = 128'h155e_340e_db25_b922_9bb1_5a2d_dceb_8029;

        #200;
        key = 128'hb657_f9e5_71d4_0704_b4e9_1b53_13f4_a9da;
        state = 128'h4934_262d_196e_6d95_6fd7_24c0_f7e3_33a3;

        #200;
        key = 128'h7b42_0f25_6a13_b59a_7148_c7d2_cae7_8a5d;
        state = 128'h91c4_016f_d255_db85_f09c_7747_43aa_7299;

        #200;
        key = 128'hfc66_1249_145c_2df6_168d_14c7_3b6f_eb5e;
        state = 128'he9f9_790e_aacb_6329_af89_2711_2cb5_f838;

        #200;
        key = 128'h3eec_7df8_495e_3303_837f_9021_460a_4987;
        state = 128'h1fa5_4714_0d29_5826_f3a5_963a_4bd3_171b;

        #200;
        key = 128'hf398_55fb_f7b0_f123_bbe1_ef1b_feee_cef2;
        state = 128'h1389_81d0_a01c_5999_528d_6330_3cdf_45d5;

        #200;
        key = 128'hcdb3_0d5a_0c2b_d220_cd38_2686_7bb8_afbd;
        state = 128'h886b_0e71_9359_37ad_cc23_492d_bccf_71d5;

        #200;
        key = 128'h08a8_4196_6b01_1961_9edd_123f_8075_a752;
        state = 128'hb90e_dfbb_6ed2_8625_6323_d830_ddef_9c81;

        #200;
        key = 128'h94e3_8a97_6812_5672_0e74_392a_fd19_8b26;
        state = 128'h445a_d585_996b_52ec_d5b9_e8b9_db6c_2f57;

        #200;
        key = 128'hef4c_c833_74b0_8617_02f1_e0fd_d918_d329;
        state = 128'hd2e8_a7d2_7102_c20a_1729_1e05_58c2_4d58;

        #200;
        key = 128'hc33b_73b0_c4d5_7ab2_2d01_0c85_95d5_db06;
        state = 128'hfd37_0812_097b_6aaa_6440_cb0f_18a1_e80f;

        #200;
        key = 128'he10f_f486_44fd_71d9_01eb_6f73_f293_da3e;
        state = 128'h6e03_43ef_50fb_ada7_f346_30db_f3c4_598c;

        #200;
        key = 128'h8028_ab7b_e303_76af_1393_0077_5ca0_c74e;
        state = 128'h7b88_dc18_ab8e_bf9c_66e8_b6fa_c971_b026;

        #200;
        key = 128'h3784_27bc_63c0_e84f_7394_afcd_53cb_348f;
        state = 128'hb69a_9113_9564_0865_b263_6b91_71ce_c89b;

        #200;
        key = 128'h9d09_8308_9b9d_0add_2a52_25f2_5b13_2d00;
        state = 128'h404b_ae61_3822_ef10_7bd3_818c_e6bf_67dc;

        #200;
        key = 128'h19ee_aa65_e1d6_bb4f_7d11_3f39_a021_dbd3;
        state = 128'h5065_b808_528b_9b48_4595_ecbe_ded2_bda7;

        #200;
        key = 128'h6588_4bd4_1f4c_83a9_da28_f173_6e4d_60c0;
        state = 128'he66c_2553_6080_3f6a_6379_48ae_f932_ac7f;

        #200;
        key = 128'h0440_14af_d9d5_4c2c_6679_30e3_7539_4805;
        state = 128'h7ed5_7489_135f_84fb_2b6e_e2f2_1f81_3832;

        #200;
        key = 128'hcb9c_d886_5ad8_4339_0f29_4256_6732_4a8e;
        state = 128'haecb_e5d3_f581_caa5_3f99_dc44_44b3_82a6;

        #200;
        key = 128'h8052_e7c5_8536_5d96_1f24_9f5e_6503_8057;
        state = 128'h390a_8eba_79f6_429b_e170_1430_14c7_3dc9;

        #200;
        key = 128'hd8f8_271e_41d7_e512_72f0_1b06_f0d7_1d5a;
        state = 128'h6c83_8f3e_8361_30f3_3bdb_ff78_4768_e50a;

        #200;
        key = 128'h9275_a88f_a1d0_57cd_41a9_42c7_164d_a47f;
        state = 128'hf3fb_3465_4f29_53cc_9594_26be_beeb_53c9;

        #200;
        key = 128'hdf52_7d63_dd82_d32f_c4e2_b1d5_ab73_eeca;
        state = 128'h45e5_ad3e_8631_06f7_b902_e36a_5879_92cb;

        #200;
        key = 128'h9e9c_a73f_2a3f_ffd2_967e_79a3_1129_f269;
        state = 128'h492d_5d03_723e_1be7_7a53_16d2_9790_4b6d;

        #200;
        key = 128'h60eb_f51a_4d2b_28db_7acc_bc74_669f_56bd;
        state = 128'h82e7_7322_bd19_00a1_205f_e4bc_903d_c359;

        #200;
        key = 128'hb133_904e_2af3_8f3c_9e14_c95a_003c_10f0;
        state = 128'h99b5_0e3b_7455_dec7_2531_36ec_b5be_46e3;

        #200;
        key = 128'hf422_812e_a619_d917_cfbb_1263_492b_0ad9;
        state = 128'h8c26_3323_7d8c_869a_26f9_a48d_4b35_9a49;

        #200;
        key = 128'hd68c_e67a_39e6_8b1b_b86d_51f1_cd36_02ff;
        state = 128'hb77a_45dc_f5ea_5b5d_4154_2f58_5e83_3a6a;

        #200;
        key = 128'h23c4_974f_c00e_88ee_968e_4747_aedd_d0cc;
        state = 128'h56ee_cd68_109a_e80a_1352_c56f_52ab_e932;

        #200;
        key = 128'h204f_6f27_58ce_bdaa_5678_9b0c_0302_3065;
        state = 128'ha2d5_7f1a_0ca5_bf0f_f0cc_6947_6e5c_272e;

        #200;
        key = 128'h599c_7260_0cfd_c9c0_b908_4e3c_c9a8_754c;
        state = 128'h6281_c5e4_840e_e7e3_8ffb_490b_ce2b_e068;

        #200;
        key = 128'he959_c96f_06bc_1beb_df6e_4e19_2d8b_26f1;
        state = 128'h99e6_550e_425e_0061_7aea_afe6_4cb2_78ef;

        #200;
        key = 128'h470a_959d_2b9b_7a5b_20c9_8d49_c572_a4ef;
        state = 128'hebe2_a742_15ae_5272_9eef_0443_5d42_11ae;

        #200;
        key = 128'h95e1_8ca1_3767_7b0c_07b7_58e1_7868_c12b;
        state = 128'h0977_bb29_6894_a5b6_3c7e_b5f1_dea8_34d4;

        #200;
        key = 128'h6613_f8c2_787d_5360_5af7_892a_0372_4f33;
        state = 128'h02ef_95d2_5439_ab40_b2eb_0c6c_5c3c_58d9;

        #200;
        key = 128'h9873_6518_74a0_fcda_8745_9201_d3b0_b2ed;
        state = 128'hc3fe_5de1_71e4_4b35_884f_800e_8e54_15f4;

        #200;
        key = 128'h868b_6087_416f_905c_4c39_cdc6_e40d_b911;
        state = 128'h7f81_a4f7_7d69_320b_bed1_dbcd_6ea7_f364;

        #200;
        key = 128'he2dc_8c65_057c_8da5_076a_8975_2b3d_e598;
        state = 128'h8e7e_49bc_bf0d_e1ec_ea29_6509_aae5_f832;

        #200;
        key = 128'h87c5_f6dd_24fe_b174_e729_51d4_61cf_bf03;
        state = 128'h82df_b03d_ab8c_7183_3572_9132_1ec5_d957;

        #200;
        key = 128'h4df6_e6c5_6b43_efe7_dfe5_fe4a_1ead_992e;
        state = 128'h42b8_19b3_7e03_111b_87fb_7e8f_773a_b0e3;

        #200;
        key = 128'h46d2_7156_99df_edcf_f53b_a539_048e_f845;
        state = 128'hae91_0fc0_0e8c_44e3_e08c_bf19_184e_703f;

        #200;
        key = 128'h45e8_6be7_63ff_ee6d_cc61_57a7_5631_0c7c;
        state = 128'h85bd_2c07_6c41_8bd2_0f6f_2d11_24bf_a824;

        #200;
        key = 128'h8c4f_ea1b_fae5_8b2e_f7e8_be35_36ec_c92b;
        state = 128'h1285_d732_a453_a58c_da3c_6be4_5542_ef05;

        #200;
        key = 128'h78f7_fb44_b498_705c_1bab_42d2_00d0_3e80;
        state = 128'h59db_659c_2621_dff4_11d9_09af_ed81_7980;

        #200;
        key = 128'h22b5_950a_23f5_f69e_4868_4ca7_4ab4_cc13;
        state = 128'hf0da_9a26_dd39_9298_a2ea_91d0_7542_fa7d;

        #200;
        key = 128'h3367_8285_09de_33ce_f5d7_9902_be86_9a8b;
        state = 128'h9f17_7987_9aa4_215f_be76_8740_a636_74e1;

        #200;
        key = 128'hc4c3_7861_ab50_1fb7_fc25_fa52_c2f8_7818;
        state = 128'h0b44_6d32_dcdf_b76d_4f14_6cc3_51b3_33ff;

        #200;
        key = 128'hbbe0_c401_7ad6_27b4_b591_f342_1b00_10fc;
        state = 128'h820d_e79e_1d3e_a8d9_0a9b_1a20_7976_786b;

        #200;
        key = 128'ha7ec_415f_f27b_5a9c_d3a2_f5bc_2c4f_7536;
        state = 128'h410d_051e_f7ff_4749_b4d0_ae24_2da7_38a8;

        #200;
        key = 128'hbf7b_d027_f910_7a66_67cc_71af_8339_4fd7;
        state = 128'hd206_9d8e_a893_8d7a_a32c_2fa7_2573_c46f;

        #200;
        key = 128'h9903_5268_1fcf_f694_5246_6095_0f4d_82a3;
        state = 128'hf1ca_0ca1_4ad6_9d75_b845_bc38_1b0c_4c30;

        #200;
        key = 128'hd46e_5db7_fc55_6c4a_de1d_e028_7e7a_df1b;
        state = 128'h108a_6a9c_8894_dd98_3d02_6792_e94a_2991;

        #200;
        key = 128'h5d74_e617_08b1_a8b7_0d22_75b5_5e8d_9c01;
        state = 128'h0739_433c_eb56_d058_58bc_5746_1cff_eb75;

        #200;
        key = 128'h7712_b165_e5e6_9006_1816_1d1f_c318_aaab;
        state = 128'h9e25_f3cf_ac37_0d80_a6fb_dcfa_8520_7ac1;

        #200;
        key = 128'h2353_c83a_e50e_e1a5_a3ab_93bc_9847_a979;
        state = 128'h2afe_2a00_3f0b_4006_80c9_136c_9160_bcec;

        #200;
        key = 128'h3c8a_35f1_f3d4_e43a_4305_575e_bec8_c208;
        state = 128'h45c7_163d_5a30_6766_1cc1_2f70_d542_dafc;

        #200;
        key = 128'h8e43_f572_50e5_4dc0_540d_75bb_8822_8a28;
        state = 128'hf5a3_f6fc_d68d_d217_98f3_1ffc_a578_1443;

        #200;
        key = 128'hdf04_469f_6ae1_d668_4c6b_e434_6791_6769;
        state = 128'hf26b_134d_6aa0_1f8a_e84d_67ac_6874_58e4;

        #200;
        key = 128'h3814_6fca_5791_2e59_96f8_b921_fd37_3a49;
        state = 128'hfe39_01c0_a5f9_beb9_ee2d_bfa8_b0c6_d5e1;

        #200;
        key = 128'h63f3_7d2b_f1fe_ae2f_9efd_fbac_5fea_6dc8;
        state = 128'hcb9b_d58e_04f8_6f04_b4cc_c778_d7a9_4a7a;

        #200;
        key = 128'ha80f_8c5d_f827_9a01_6dbd_8bd2_755e_d091;
        state = 128'h77ec_4b4e_71a8_9465_407e_566b_b13b_3edd;

        #200;
        key = 128'h5527_2bbd_d399_0ada_3836_874a_4f9f_a2d1;
        state = 128'h3f07_5531_46e7_f7bf_bf6d_c36c_4cc2_4d14;

        #200;
        key = 128'h52fc_f449_6b96_484a_c71b_29c7_aee7_5798;
        state = 128'hdd53_f139_150b_9074_2411_6d03_d36f_427c;

        #200;
        key = 128'hc472_7562_a754_2d3d_fa84_ed77_a23b_01c4;
        state = 128'hf989_48a5_9d31_f993_15ea_0c6e_b9cc_09bb;

        #200;
        key = 128'hbbb0_3417_bc20_daa2_3c35_655a_aab8_e02b;
        state = 128'hce4e_e229_441f_3381_3569_c792_b955_25d2;

        #200;
        key = 128'h9639_2976_fe90_cc10_81fe_2404_695f_456a;
        state = 128'h0a06_b7c6_c804_9b3a_1609_be3e_a746_c1c6;

        #200;
        key = 128'h6984_af31_02b9_2184_222c_af4a_67c0_93b9;
        state = 128'h0dba_5c79_3314_ed74_228e_5f31_a230_3d6e;

        #200;
        key = 128'h5564_4d59_00a2_9ac2_d827_5344_a953_1df8;
        state = 128'h48cf_f75d_008f_79ec_9d83_8a35_2674_eae3;

        #200;
        key = 128'h0a94_51c2_a5fc_0a29_b4c5_b115_d7a8_83ba;
        state = 128'h2878_6b65_baef_5ad9_d3bd_5959_0e8a_08c4;

        #200;
        key = 128'ha8d7_c82f_4c37_efbe_45c4_c833_18b1_6ee8;
        state = 128'h5679_3fdd_88a8_0aca_5536_c69a_319c_cf38;

        #200;
        key = 128'hcf17_74ee_4b54_0d7b_ac95_6f7e_477b_026f;
        state = 128'h2e80_bfaf_0a62_f13d_2951_4e3f_cf57_a261;

        #200;
        key = 128'heb07_dd13_a739_2c8d_971d_a0c2_c02e_448b;
        state = 128'h2134_9ba1_fdb6_abe9_8bab_c286_a033_a809;

        #200;
        key = 128'h6a93_82af_fb63_2bbb_83a4_4892_dc87_4306;
        state = 128'hf878_0a58_4c82_45d7_6a21_9d2b_a4e5_b550;

        #200;
        key = 128'hfd23_8bbc_6ef0_55e8_5bf4_29b2_6d00_2c05;
        state = 128'h36ca_6c0c_3bd9_6146_8d9e_6e75_a359_766f;

        #200;
        key = 128'hc97d_81c6_2475_667c_bae0_1e35_7384_ee64;
        state = 128'hdba4_3d2f_d80c_f286_5dd7_0836_2d68_68db;

        #200;
        key = 128'hde1d_74e2_4368_d40b_3aa4_c10f_eaa6_5004;
        state = 128'h98a0_a901_1371_bf62_70a3_5c55_d497_8b57;

        #200;
        key = 128'hab03_4bd9_ba33_b5d1_fdac_076f_71a5_3304;
        state = 128'h0a8a_66ab_2406_750f_f552_7e6b_23cf_02df;

        #200;
        key = 128'h0e5e_fd05_3518_e6c8_cfb7_5795_598d_8cce;
        state = 128'h4e4d_40ea_7531_54b2_3ec7_79ff_b835_7f50;

        #200;
        key = 128'hced2_f399_d0b3_61df_dabe_41b7_bb8a_6de0;
        state = 128'h2ac0_64e1_35fe_0894_dbb3_f8fd_ab50_132f;

        #200;
        key = 128'hf5ce_e03a_2eda_ec27_be79_9084_c071_81ae;
        state = 128'hed19_b1ae_dc1b_3503_5476_39fe_0c0d_0032;

        #200;
        key = 128'h1a3c_5f5e_52ce_c566_d526_e23e_7d5f_bce8;
        state = 128'h740d_4c8f_93a8_28e4_83d4_70f5_58dd_4ccc;

        #200;
        key = 128'h5836_ab51_03fa_e305_86a5_2667_6736_f6a5;
        state = 128'h1eb9_0d7a_3184_915e_51fd_e08b_06c6_295f;

        #200;
        key = 128'h1f57_9a34_fb2f_b199_18bb_cd3e_2c8b_0cb5;
        state = 128'h13b3_2737_1ec0_9ec6_1081_e7e6_5591_483e;

        #200;
        key = 128'h9531_c962_9c5a_430a_dd17_d1a3_6ab1_1c89;
        state = 128'heee8_866a_b370_8891_06e5_2eb0_3ec3_351d;

        #200;
        key = 128'h5bb1_f0e6_c028_7cc9_b956_383f_04d1_5d95;
        state = 128'hfb4b_e976_7827_438b_f5f8_48e4_0694_fb79;

        #200;
        key = 128'hf0b0_5dcc_7ac7_f946_146a_ab28_2353_76bc;
        state = 128'h8515_bdf5_7b80_6c20_1c50_e3dd_2d58_3bf2;

        #200;
        key = 128'h68a7_f251_d4b1_5e10_4d84_91f3_210e_bf76;
        state = 128'h5b95_790b_ed20_3dd6_2b9d_5ab3_b92d_6f14;

        #200;
        key = 128'h7b34_a61b_445f_7299_96ad_4f83_5c60_261a;
        state = 128'hfc5c_096a_9f1d_23f0_54ee_c843_bbbc_c419;

        #200;
        key = 128'h4775_4875_290d_90b0_60e1_a1d6_1b36_fae3;
        state = 128'hb5aa_951f_4e3c_579c_b973_8edf_9ec6_d622;

        #200;
        key = 128'hc9be_4631_eab4_3f69_4eb3_0a67_8daf_eec8;
        state = 128'hf84d_ab27_67ea_bd72_2c41_5281_936c_298d;

        #200;
        key = 128'ha2ff_dff1_0821_300c_53ab_68bc_ac0f_d1c8;
        state = 128'h3582_9198_c3ca_1a5f_bb35_6b9f_cd04_2023;

        #200;
        key = 128'h9575_cb53_c686_d419_fc46_a417_158e_ebb8;
        state = 128'h8ba5_0d88_59a9_6cb2_4d0c_937d_fa3b_7c5d;

        #200;
        key = 128'hf553_627c_167d_3aa6_541c_4fa2_380d_9108;
        state = 128'hf770_413b_a2ad_7053_7f4c_0bad_26fb_a3ad;

        #200;
        key = 128'h86d5_7b7c_58ac_ac62_82a3_bd2c_2868_f870;
        state = 128'h7030_f3e2_2ab2_dd15_ac23_b97d_4b30_ff2c;

        #200;
        key = 128'h6c3e_fa24_db93_b18a_4dc5_7b9a_3b24_1f88;
        state = 128'h100a_5dd2_5639_a407_326c_fb9e_5917_9c0a;

        #200;
        key = 128'hb305_b46f_ca9d_0e0f_5d15_b490_0c16_ef68;
        state = 128'hc2cf_84f6_ea6b_b185_1c20_342a_780f_6d8c;

        #200;
        key = 128'h58ee_dc4d_e9fe_bc93_2974_2b50_fbeb_01bb;
        state = 128'hc544_bafa_8a6a_5ebd_056a_7e89_4f66_929a;

        #200;
        key = 128'h3016_a340_2f4a_720b_9760_1824_b024_b7f9;
        state = 128'h48c6_ed93_8353_7ddd_89fe_c2a5_2b74_f622;

        #200;
        key = 128'h8c49_9acb_a7d9_2d82_ff74_487a_2c75_6c29;
        state = 128'h35dd_915c_1863_d545_0df0_7375_8979_c3cb;

        #200;
        key = 128'h0071_52f9_578b_5e9e_8c92_f742_a007_a02a;
        state = 128'h6098_9e2b_1cc1_b1a0_cf22_85a4_c704_00a6;

        #200;
        key = 128'hada5_cc4e_0495_fd27_4039_fcb7_3610_14f5;
        state = 128'h50e3_0bd6_44c4_fbc4_33b2_dc53_59d7_bbf1;

        #200;
        key = 128'h8861_b8b6_aa9c_7583_8995_7f9c_a9c8_10ac;
        state = 128'hc7c7_989c_4f01_a6bb_8f4f_6b9f_7ae3_eb33;

        #200;
        key = 128'h9613_c49c_1a68_6b34_5f66_db19_d429_80cb;
        state = 128'hb1f1_2ede_a078_84b1_f1ab_5830_e892_064f;

        #200;
        key = 128'h48bd_b598_d30a_67cf_af50_b59c_1888_ff92;
        state = 128'hf08e_127a_4299_ef9d_327a_9214_b1ed_f7f0;

        #200;
        key = 128'h47e5_aa58_427e_b1f3_3009_3f06_1b19_3b35;
        state = 128'h5147_09c4_ccb3_768d_368b_86d3_dae5_238a;

        #200;
        key = 128'hb629_e920_a793_c6bd_07be_101e_1f82_98f7;
        state = 128'ha829_6ef6_d494_a8ae_4bb0_63b3_f0fd_6aa1;

        #200;
        key = 128'hf0e2_1095_e3a7_e8c7_3a4a_a2f0_2343_9e5a;
        state = 128'hf35e_18d0_6ec1_ca5e_cd60_5c5d_5acf_e0ca;

        #200;
        key = 128'h7151_6958_9936_5f73_e9c5_5660_de4e_4169;
        state = 128'hfdbc_4156_4060_3e13_9981_86f0_ac9b_1667;

        #200;
        key = 128'h0a56_b7eb_75c5_5d58_2913_2626_bd57_598b;
        state = 128'h2d40_046e_40fe_de10_93f4_412a_fb80_7cde;

        #200;
        key = 128'ha2e7_8655_6b24_da32_d968_2cab_2ec8_fc77;
        state = 128'h4bcb_2866_de74_413f_b337_5179_5d40_0698;

        #200;
        key = 128'hd074_ffdc_b332_72e5_1792_a16a_e264_8243;
        state = 128'h49b9_f563_f495_6b08_cfc9_c948_b5e4_7633;

        #200;
        key = 128'h337b_3ab1_620d_e860_d89a_18cc_a466_d599;
        state = 128'he42f_7845_afa3_f0da_b022_a575_c800_b264;

        #200;
        key = 128'hd64f_7172_dff9_e188_841b_35aa_1a9f_ebf5;
        state = 128'hb6b1_c8db_03e6_2013_f093_41b7_7da5_1b1c;

        #200;
        key = 128'h8f16_1641_0c99_3469_63f4_95cd_3a5e_bb43;
        state = 128'h46e6_d039_d879_88d9_06b2_bc5b_60b2_6df5;

        #200;
        key = 128'h871e_1d01_f186_9b10_3014_42da_a8f6_4029;
        state = 128'h7aed_c7ea_3443_b3a8_1fd9_ad24_15ff_5c77;

        #200;
        key = 128'habc1_86ac_4e49_7b13_7b93_02c7_143f_f5c5;
        state = 128'hd305_7494_209c_5cb6_1d14_c08a_9d3b_16aa;

        #200;
        key = 128'h8f0e_4298_3ccb_7c78_5b44_fc06_5bb4_a7f9;
        state = 128'hf077_a636_e9fe_bbd0_f6b2_c76f_f440_7bd6;

        #200;
        key = 128'h7525_e51e_b075_eff6_d182_45bf_e560_d1e5;
        state = 128'hc6d1_a85f_6dbe_a366_5c0a_52ac_8334_052c;

        #200;
        key = 128'h8414_8695_e294_38c0_5172_274b_8586_4245;
        state = 128'h8096_9ddc_3504_50d5_a233_e598_7d22_fdd8;

        #200;
        key = 128'h5bda_71c5_05a2_14e0_18d4_ec6e_a15a_48c1;
        state = 128'hb5b8_3fef_d315_d647_4c01_6d11_2398_28d8;

        #200;
        key = 128'h8cc2_63b5_89bd_6f26_0281_3fca_2830_4af7;
        state = 128'hc7d2_d26e_90ac_35b4_3814_7317_b452_d20a;

        #200;
        key = 128'h0c6b_aa32_bc2f_c8d0_7372_d659_d432_5d8a;
        state = 128'h926c_de7d_920e_5698_198a_fe82_c384_84ca;

        #200;
        key = 128'haeab_bff2_5a43_8d4a_f348_e3a8_6a94_e726;
        state = 128'hd285_c2b1_4666_93a5_e47a_2780_2d30_af8e;

        #200;
        key = 128'h33be_dc55_e632_a887_dd69_0d65_f629_757e;
        state = 128'h56f3_cadc_5b6a_444a_196d_8b0e_2f16_d65f;

        #200;
        key = 128'h3f68_740f_1651_8f7a_b519_3805_b031_cec6;
        state = 128'h917e_b229_00f3_38e8_063f_5353_dcb2_5f19;

        #200;
        key = 128'hae4b_c575_01aa_5b0a_e7b0_2c99_f6c5_5b63;
        state = 128'hfbd9_cca1_e307_dff9_c9ff_5b4b_fbfd_c1e6;

        #200;
        key = 128'hf457_e74d_436e_4141_b132_06bd_4120_d5a7;
        state = 128'hf4a9_ba44_5fc6_380b_f606_699c_4766_6195;

        #200;
        key = 128'hdfa1_ac74_c167_e2e5_11d8_601d_d4e6_b0f8;
        state = 128'h33ea_336d_7704_2b66_c95b_ab83_1a8f_9dfa;

        #200;
        key = 128'h7be2_8b52_9257_a2cf_0b71_88dc_a855_9046;
        state = 128'h5e0e_b1ae_95fe_b19f_c521_1af7_e314_9d37;

        #200;
        key = 128'h76be_aea8_95dd_3b79_14b8_1968_0080_28ce;
        state = 128'h5542_f0c9_2d28_10a1_7eb9_b0b4_db5e_d618;

        #200;
        key = 128'hf73f_2219_2863_aa41_2de4_1416_083e_171c;
        state = 128'h3182_270a_50cc_e0bd_8f7c_c5ef_60c2_2ef8;

        #200;
        key = 128'h2e80_5ed1_c22b_d1f4_c1fe_e3e6_f53a_222c;
        state = 128'hd56c_4701_799e_3024_effc_e481_1c25_48d6;

        #200;
        key = 128'h182d_7198_a396_1270_8a5c_774f_40c9_8c1f;
        state = 128'hc057_8a4a_f06b_10ae_51b7_98e1_26db_caf1;

        #200;
        key = 128'heec8_dac7_8c49_a29a_6998_75a8_114b_f56d;
        state = 128'h7831_8c28_72c2_e9f4_5fa1_92e2_ae9c_c25f;

        #200;
        key = 128'h55a9_1756_b904_cb1b_6e40_5e59_624b_6b65;
        state = 128'h32f8_74b0_28ae_7089_c943_9bad_5787_7cf3;

        #200;
        key = 128'he941_4115_31e1_1e13_45fa_62cd_22bd_7927;
        state = 128'hedba_1a0e_4d6e_41f1_d238_af91_ff41_e2c3;

        #200;
        key = 128'h0e7c_a051_ab1e_8610_1fb8_d34e_ccf1_151a;
        state = 128'hc2c9_e45a_d063_438e_e56e_11b9_6b84_30de;

        #200;
        key = 128'hc513_8af0_9df6_9b7e_0c90_5bef_0c49_6685;
        state = 128'h082c_e221_33b8_8254_78d0_b8f7_5e66_658f;

        #200;
        key = 128'h2700_03cc_4ac5_dc4c_2741_8c21_b931_8aa0;
        state = 128'h8ec9_2011_95dd_584d_69be_50a7_0177_96ce;

        #200;
        key = 128'ha6ec_c07a_84ec_5472_e0d6_f771_938b_6aa1;
        state = 128'hc311_1df1_0ed8_e93d_bf9e_27f2_4bc7_c29d;

        #200;
        key = 128'h004f_c93d_89c5_7b8c_2d5f_0338_c60a_a7b8;
        state = 128'hbdca_630e_06e5_5844_68dc_94f1_da2b_2885;

        #200;
        key = 128'h08aa_d972_d7f1_b341_a039_6347_5eee_bc2b;
        state = 128'h0ee2_e866_ae43_e3ff_7e96_802b_382d_1624;

        #200;
        key = 128'h1c6f_16f1_6e28_0adf_e1f3_1543_e6bf_45e6;
        state = 128'h394d_771c_0283_1d48_aa0b_1311_d961_b32b;

        #200;
        key = 128'h9af0_9217_1d71_7f99_1857_4527_d41c_dbb8;
        state = 128'ha944_8046_8dff_faf4_8104_3a78_1f3f_8313;

        #200;
        key = 128'hb80c_5a2e_88b3_df04_b2c7_9fbc_ade2_d1d9;
        state = 128'h210b_299d_c159_e107_1837_cb64_884a_ac82;

        #200;
        key = 128'hdd70_5997_07de_65a9_1987_3b6a_8c1b_5cb5;
        state = 128'h332a_1c00_058c_2da9_ba18_66f7_17e4_f3e1;

        #200;
        key = 128'h7dbf_7097_7fab_66e0_0c1c_2a6e_14f2_e6c1;
        state = 128'h4e09_225b_95fb_7fce_1ae4_ede0_9bdb_42af;

        #200;
        key = 128'h4c4e_234d_70a8_2c05_fc15_7956_0536_264c;
        state = 128'h0b8c_f45f_fd55_0313_1a87_ec09_dc9f_74db;

        #200;
        key = 128'h87b1_88fb_d00d_677c_1dca_8cb0_02fc_2ede;
        state = 128'hfad3_5b76_a5d7_956a_4021_6a52_cd9b_239a;

        #200;
        key = 128'h0cc1_508b_e135_0237_8db4_3daa_d79d_8217;
        state = 128'h2362_b86d_2893_0801_40e9_1712_abfa_6756;

        #200;
        key = 128'h9f24_6036_6c8c_a2c9_6d40_3004_3834_d72c;
        state = 128'hbd61_436d_e479_2d12_c775_789f_7be5_1515;

        #200;
        key = 128'h60aa_61b9_fedb_4d42_a830_a692_658d_ef00;
        state = 128'h2e6a_6c05_b92a_b50f_4465_aa90_00ba_71ba;

        #200;
        key = 128'h5cac_5d4c_841b_93e0_55fa_3a47_74cb_acfb;
        state = 128'hfc5a_b3f6_5159_ca55_2e97_aadc_c2ad_0566;

        #200;
        key = 128'h010f_4908_d362_a7ee_5534_af20_6152_cb11;
        state = 128'hd798_9a81_7d36_cd31_444c_b680_69f3_4961;

        #200;
        key = 128'h15c2_aa4d_36db_852a_e559_30a6_baa3_cdec;
        state = 128'h7517_ac49_7644_1000_a6ae_1d2e_c839_64a9;

        #200;
        key = 128'h5fc8_c0e2_8212_8680_8a56_8e33_60d3_7320;
        state = 128'h0817_f38d_d79b_0511_1f01_1dfd_3b44_6541;

        #200;
        key = 128'h8cde_e267_e9f8_34dc_4eea_5c19_70c4_c752;
        state = 128'h049a_71b9_4003_e2f9_386d_b2d7_af96_62ed;

        #200;
        key = 128'h6b4b_ae99_2333_096c_4699_b249_f533_e659;
        state = 128'h2791_b94f_2287_a3c1_a51f_ab2f_546e_fc3e;

        #200;
        key = 128'hb26f_a4be_048b_ba9d_9163_a3d5_269c_b948;
        state = 128'h3551_aff1_a9e0_ea3e_1ae1_e061_ca52_1ff9;

        #200;
        key = 128'ha7b7_fa3d_f17b_1b04_8bdc_bbff_3972_2814;
        state = 128'h9d12_99a9_7a01_71f3_f608_385a_dc76_f497;

        #200;
        key = 128'h13ff_1cd8_b124_f2fe_0247_7994_b025_1a85;
        state = 128'hb8eb_01b5_fb50_f1a2_1429_86ca_3584_11fc;

        #200;
        key = 128'h71b8_7d31_346f_6605_a5d5_3b08_89e9_b304;
        state = 128'he639_56b2_b1c1_0ec0_df82_89de_4cf8_58ad;

        #200;
        key = 128'h0bd0_876f_2bfb_1615_1814_4f7f_16e1_31c0;
        state = 128'hc7cc_2d19_852b_f18d_8566_920a_3a89_95f9;

        #200;
        key = 128'ha324_7a27_e76d_94be_d29d_b58c_7e4a_ffbd;
        state = 128'hb00e_df7c_e294_eb31_ced1_b841_c8c7_baa3;

        #200;
        key = 128'h23fc_17ae_310d_3e28_1701_5b65_d667_1715;
        state = 128'h892b_eedb_2f47_909a_183b_f6c8_35db_9b45;

        #200;
        key = 128'hac9d_e7f6_1f30_2382_9e3c_0001_1d64_f918;
        state = 128'h763b_f455_d2a6_af29_258a_28a0_8123_c62f;

        #200;
        key = 128'hc4e8_cc3f_ad7a_b944_44bd_7275_96ed_742c;
        state = 128'hd863_1e3c_9a08_e1c0_c712_407f_1a1f_b5f0;

        #200;
        key = 128'h1789_e5ff_e83d_c942_6853_605a_bed6_1836;
        state = 128'hb2ac_ba75_28c4_36b6_4714_9538_5582_eb2d;

        #200;
        key = 128'h5c73_a068_147e_4742_b1dd_2dc5_30ac_85db;
        state = 128'hf2d5_a96d_ee5e_8f7b_5fec_5aa8_8a43_f6af;

        #200;
        key = 128'ha1b5_d3e6_61a1_5fed_2583_cabe_d401_4ad5;
        state = 128'hda60_930b_5c3a_9117_ee83_c1a8_f9e8_5d06;

        #200;
        key = 128'hefaa_2c0f_98ab_fb2c_a10d_fa8d_5efe_af76;
        state = 128'h584d_24bc_d88d_7b59_aa51_7e19_3feb_71d0;

        #200;
        key = 128'h6796_8697_957a_4578_3f3a_1d01_86e1_8b45;
        state = 128'had85_06d6_6101_a84c_ecfa_e209_326f_7806;

        #200;
        key = 128'ha236_3328_5c4f_fc86_09dc_0e02_e62d_1557;
        state = 128'h2c27_fcd3_8b22_8b97_7c01_6b0b_28dd_e569;

        #200;
        key = 128'he373_8de7_ee79_e66c_64c5_0c24_a779_0edb;
        state = 128'h6c7c_ef08_f098_7ce1_e1e4_3f81_404c_b27c;

        #200;
        key = 128'h3ad4_21a5_2af0_2a0a_a123_84c8_8e74_c902;
        state = 128'h1eb7_cb51_4e76_0b83_5d2e_afc4_ea87_cbef;

        #200;
        key = 128'h6d5e_7e34_e415_16c7_0ff5_eaea_b5bd_e461;
        state = 128'h8854_22e1_b94f_0b2c_7e78_80b8_fed2_9ad7;

        #200;
        key = 128'h43e4_7a42_08c0_e6e8_8734_1e2a_fb16_34ee;
        state = 128'h4498_f078_a613_3695_faac_a1b6_3e52_fb5f;

        #200;
        key = 128'h2e24_e3ea_40b2_f8d0_3609_e6d1_3116_da3e;
        state = 128'h529c_cc2f_13ab_92e4_b633_ef4c_fcca_466c;

        #200;
        key = 128'h2a85_12f9_1164_469b_4b02_3c28_bcdf_3463;
        state = 128'hbb7a_609e_07d7_d724_fe0c_6e9d_0990_196e;

        #200;
        key = 128'h5309_f150_35d9_baf3_9382_eac0_232a_2c46;
        state = 128'h4352_1529_7841_7db9_053a_c435_8e4b_696e;

        #200;
        key = 128'hc866_e602_c2ff_e3ef_89c7_1226_833f_ed8e;
        state = 128'hd5fe_7a3b_e869_f91d_aa17_22d6_6a5d_dc11;

        #200;
        key = 128'h5005_d126_9d45_96f2_bdf3_31f5_930f_8674;
        state = 128'hceb8_7d00_5e7c_cfca_9abe_5e0b_b45e_dd30;

        #200;
        key = 128'hdd28_6605_b5ff_56c2_b030_16bd_2fb3_9443;
        state = 128'hd058_6037_6757_1d1e_35eb_3e0a_d205_2048;

        #200;
        key = 128'ha9f7_2038_dbc9_de44_ce96_1dc3_ebfe_76c3;
        state = 128'h3382_1de8_9fd6_22de_da20_3804_49cc_1506;

        #200;
        key = 128'h07d8_d98a_3fb6_cb26_8be0_66ea_640c_3c0e;
        state = 128'h5c03_c52e_c805_dc9d_a3d5_7074_c828_cbd7;

        #200;
        key = 128'he38e_6b1f_baa2_ce32_0d9c_8e0d_a835_3eb7;
        state = 128'h4cc3_f089_9f31_1b0e_8398_2543_ed1b_2149;

        #200;
        key = 128'h92b9_5d3d_48c1_1b27_25ae_4b09_763a_3019;
        state = 128'he29e_6d95_e52e_ef5d_a3b5_f00a_8bc7_7475;

        #200;
        key = 128'hc0bc_1752_5234_65f3_817c_02b5_6b82_b3d3;
        state = 128'h9179_bda7_caa4_9ac3_4a24_1d10_a7a2_5817;

        #200;
        key = 128'h0e21_79a1_670d_aa43_109a_ec8e_0c43_bd8b;
        state = 128'h8330_a08b_9318_c872_4070_0abe_0c41_13a4;

        #200;
        key = 128'h7c7c_c975_5fa8_c183_531a_5437_d3c1_a8c0;
        state = 128'h3d85_533f_0150_e7f9_5531_4e0a_b80a_141b;

        #200;
        key = 128'h5c29_4323_2da9_2af5_1de4_3c12_b3fc_f400;
        state = 128'h2bf5_4dd6_ab80_c711_fc39_a684_5cfa_eeda;

        #200;
        key = 128'h4048_8910_2d04_8c1a_0627_2078_e82e_86a0;
        state = 128'hec8d_ceaa_c9f1_32da_27c9_b6d5_a2a6_4c3e;

        #200;
        key = 128'hcf28_eaf4_47f8_197e_7f4a_f240_acef_fa5a;
        state = 128'hec00_a23f_f9cb_4232_7afe_25ea_280a_df4e;

        #200;
        key = 128'h799e_bba3_9c0b_9362_bf0c_db9e_6002_1122;
        state = 128'h99c0_822b_44b7_c399_3f8c_6bcc_bf2a_a36b;

        #200;
        key = 128'hb6ff_c93a_8448_5f63_4bfd_933c_a632_0c7d;
        state = 128'h1ba7_bad3_d8dc_9048_f66d_1b1b_92a9_1f6d;

        #200;
        key = 128'h48fe_5f9d_1e05_0e08_a682_25ef_6601_6b61;
        state = 128'h8e12_3f5f_15b4_3653_b015_b75b_4be7_ef3b;

        #200;
        key = 128'hdd28_6dba_d3eb_b8ef_b10f_2b80_5303_8f98;
        state = 128'h0886_c5a1_e2c4_8e8a_201c_bead_a347_404d;

        #200;
        key = 128'h0dc9_ae52_4057_8b03_2632_a2ff_c8b5_f2c3;
        state = 128'h56ff_3345_2156_0222_47f5_c2b0_00d2_0f11;

        #200;
        key = 128'h6e18_c54f_fb22_f893_53cc_7a4d_b26a_581e;
        state = 128'h336e_153c_cf20_9db0_a897_9bf1_510e_3846;

        #200;
        key = 128'h7584_ca3f_5fef_4700_362c_d692_78c1_345e;
        state = 128'h9e56_4fb0_ed11_0a7f_e4e6_c78f_1287_7986;

        #200;
        key = 128'h7e79_f47a_7fb6_afcf_38a2_f5a4_f980_eb0a;
        state = 128'hb944_a077_67c1_a820_1605_e7de_0c22_2329;

        #200;
        key = 128'h38d9_a830_730e_bf66_a61f_d044_0233_7b32;
        state = 128'hff41_5e76_1b06_1473_94a2_6dfc_0099_60bd;

        #200;
        key = 128'h5887_8af5_744f_c1b6_c7ed_c5df_8cf3_0329;
        state = 128'h85e6_333f_56f6_31f9_7847_19b0_3029_f646;

        #200;
        key = 128'h93f6_a936_24e3_c3cb_c44e_7816_2f40_ac08;
        state = 128'h06e8_3d4d_3288_06a3_2784_7ac4_003a_4fd8;

        #200;
        key = 128'h878a_d623_35f8_34b8_6466_2098_b36d_5dd5;
        state = 128'h2560_e440_4262_11dc_fb53_b469_3963_d5c1;

        #200;
        key = 128'hca27_4613_5add_c936_8f3f_e85e_1b57_6527;
        state = 128'h39f6_4461_182f_60ef_9e79_b6be_0fe6_27fe;

        #200;
        key = 128'hfa3c_10fe_c4b8_84c0_6e68_c3eb_f853_9b63;
        state = 128'hb2e9_fda9_df9d_f7b2_d749_a9a2_a7b3_1f3e;

        #200;
        key = 128'h1645_4bfa_e89d_20c9_ee7c_b069_47b1_5c33;
        state = 128'h24b7_3aae_24ea_3e98_8bca_659f_e243_0552;

        #200;
        key = 128'he83b_489d_74a5_cc36_6292_0edd_28f0_23b4;
        state = 128'hd0cd_1d98_36d1_4cb5_5700_efca_c907_7959;

        #200;
        key = 128'hb820_91b9_8f13_b652_5c4a_1c19_08f9_2fbf;
        state = 128'h90fb_ba86_10ad_a243_7712_e6e8_6638_5948;

        #200;
        key = 128'h828b_5efa_1bef_f9df_716d_e917_e58b_321c;
        state = 128'he451_79a9_805c_d0ee_c109_d460_b40d_f967;

        #200;
        key = 128'h3bfe_2f47_f078_c361_337e_7bc3_1425_e4f3;
        state = 128'h2a52_b9c5_a253_593a_19fc_2fa4_c889_e2bb;

        #200;
        key = 128'h5817_7270_54d5_c1b1_5e58_d2ff_2b49_b989;
        state = 128'hf331_4549_a777_fa1d_b970_6fb8_c256_fb27;

        #200;
        key = 128'hb276_5256_3c0d_76ea_e8b4_a0d7_d800_8009;
        state = 128'h00c1_6f3a_2949_3617_2719_f33f_e832_2bcc;

        #200;
        key = 128'h62dd_cd49_fef9_a9c6_7d39_708e_edbf_e5cf;
        state = 128'h1214_cd5b_c4b7_0e57_5c93_e806_b640_d614;

        #200;
        key = 128'h1af4_ad44_b328_666f_c6dc_187d_8f1d_f7ae;
        state = 128'hdc7f_61a5_043e_c657_07b4_2f6b_8fda_22fc;

        #200;
        key = 128'hb6ab_bf7e_2421_e1bd_35ec_47ed_3a96_e70f;
        state = 128'h33a2_0127_6be6_e71e_98b1_62b8_e25e_b426;

        #200;
        key = 128'h98ea_e225_2902_c3ce_b630_3bf0_5b08_b6ed;
        state = 128'hd4c2_5962_ccea_6863_ef19_83d0_5709_fc04;

        #200;
        key = 128'h73e0_6bc5_073b_2381_be75_12b5_bdd8_6c33;
        state = 128'h3d7f_120a_cf08_b20b_8ecf_b8a5_0386_d389;

        #200;
        key = 128'hf7b8_8faf_82f4_8f80_8192_06aa_4d02_58f3;
        state = 128'h7c02_6992_93bd_6f82_2a15_8baf_dd3c_074d;

        #200;
        key = 128'hca9f_b537_cce7_e983_e296_ee30_7dd2_57bb;
        state = 128'hb46e_9ccf_a180_833f_0ff9_8182_7117_9220;

        #200;
        key = 128'hc20f_32ea_d14d_e23a_cd0d_81db_72b6_51dc;
        state = 128'h1dcb_9100_151a_a792_9812_c2ac_0787_07ff;

        #200;
        key = 128'h55fc_60bb_cb79_5b6c_eb9c_144c_9c1f_75a2;
        state = 128'h56c4_3de9_c46e_908c_946a_39b1_d2f1_58c9;

        #200;
        key = 128'hc9f3_947f_7a99_58fd_f66c_84b7_7426_95b6;
        state = 128'h6a13_dcc3_c98c_dba0_af5e_078d_ca79_b0a5;

        #200;
        key = 128'h87ed_056e_503a_1a1c_80dd_28b2_875c_98de;
        state = 128'h042b_2729_b3fd_4341_e150_2570_48c5_ab6b;

        #200;
        key = 128'h676f_11a0_577b_6b12_7ec7_0664_fc45_ad25;
        state = 128'h5d65_fad3_2142_9939_0f2b_42e7_b9a4_1779;

        #200;
        key = 128'h22c6_6b41_29d8_6dcb_ab29_0106_5e5d_b9da;
        state = 128'hb924_1370_fb75_062b_0bba_c4d2_31fb_86a9;

        #200;
        key = 128'h3f1c_4ff5_3ce4_988b_f899_caf8_d0f9_5890;
        state = 128'h03c9_34b0_418f_a3d9_85ae_cc19_2bb4_2001;

        #200;
        key = 128'he288_73ec_9965_7e32_beaf_d910_0689_1c54;
        state = 128'h0135_8e30_88e9_915d_0ef8_5d02_2fd8_98f5;

        #200;
        key = 128'hb965_dd24_3103_e504_4fd8_f62a_8771_a35b;
        state = 128'h78d5_c95f_2b42_24dc_e03d_6929_312f_d91f;

        #200;
        key = 128'hddc7_9b83_8f5d_d5bc_efa3_636c_de0f_6c0a;
        state = 128'h6631_14f0_c7e2_118a_0e48_9a28_8f53_3033;

        #200;
        key = 128'h5818_5a90_4524_61ad_77f9_7b33_ad41_3991;
        state = 128'h15cd_451f_e961_a55c_b0a0_5d27_48aa_c95f;

        #200;
        key = 128'hf010_9b5c_ebfa_aebe_79c4_c587_b431_08ef;
        state = 128'h7b7e_e910_5a63_1867_5096_2020_2958_6e3c;

        #200;
        key = 128'ha548_c172_4eca_4a05_d60d_477d_3a83_378c;
        state = 128'hf7c1_07e8_d7a7_6f28_6723_5488_e3d0_4e2c;

        #200;
        key = 128'hc0e3_4362_a48d_e14f_f431_69d9_eb40_c593;
        state = 128'h3256_747c_c87e_c78b_b93d_1240_31fc_09dd;

        #200;
        key = 128'h6ae8_9c4f_d38f_13dd_0672_fd1b_93d6_5ec9;
        state = 128'hb1c7_3297_4f48_9768_17ca_5d1b_16e6_a1b8;

        #200;
        key = 128'he33b_75b8_ff6a_5671_8c3c_747c_e488_83af;
        state = 128'h74b9_40e7_2c88_a2dc_367f_c928_db4b_02b9;

        #200;
        key = 128'he9e7_9ffe_8b3b_880c_366c_f582_7a10_26d6;
        state = 128'h2573_589b_ce0f_bd07_4d95_0606_bffa_9279;

        #200;
        key = 128'h4a00_e28e_2f8c_1274_7008_3c96_97e4_4174;
        state = 128'h8973_d1cd_61a7_0849_c1d4_cc85_ef7a_0168;

        #200;
        key = 128'h9599_6e73_8c11_669a_66ed_63e4_dc19_58f1;
        state = 128'h58c6_b6d9_ec07_0966_c3ec_25e7_a18f_2451;

        #200;
        key = 128'h2281_aac4_0bac_88a1_de41_be3c_cd99_f700;
        state = 128'h7b26_75c7_a031_b211_b918_2345_4aa2_425b;

        #200;
        key = 128'h9d87_be38_d151_7f85_6e48_869a_deb2_a76a;
        state = 128'h28a6_a7fc_5a8a_3655_b89e_305c_839c_ca43;

        #200;
        key = 128'ha084_2c7b_cce6_e9ce_7b71_b12b_ea2d_e047;
        state = 128'h70fd_0147_3aad_982f_e0d2_3689_4c76_40ae;

        #200;
        key = 128'h3075_bd31_483a_5d42_984f_87f0_4fbd_0e87;
        state = 128'h8fdf_704c_653b_5624_094b_1acb_2274_4627;

        #200;
        key = 128'h3478_22cc_e48d_1d3a_c141_4924_3ac2_84ac;
        state = 128'h12b2_d20e_fc4f_6231_9e15_313f_75a8_9df9;

        #200;
        key = 128'he5fa_3716_c2b1_5a25_d644_e702_9b77_f11f;
        state = 128'h711f_c98a_620a_2dc7_71a7_f197_ba3a_0b17;

        #200;
        key = 128'h4405_4a33_fe58_d64d_b784_9fce_4b53_944c;
        state = 128'h81ae_fd68_92b6_9a00_41f7_88d9_c2f3_a002;

        #200;
        key = 128'h50c4_53cc_3ffe_307c_d676_f54b_1b77_ee34;
        state = 128'h9db2_7554_4997_45a1_6e34_4238_b26d_02dd;

        #200;
        key = 128'hd727_b2bc_d3ef_ac49_8d17_fe44_8bf2_1b58;
        state = 128'hcefa_cbd3_e19b_7ebd_fed7_f4f2_0690_4af2;

        #200;
        key = 128'h629f_ddd2_3eba_e770_e1ee_6dc3_eed7_6daf;
        state = 128'h8186_915c_d7eb_e6ce_85d4_a701_64ef_8e93;

        #200;
        key = 128'h6e15_0558_0b2d_ed4f_e62f_4110_2909_2687;
        state = 128'hfc8f_0f9f_5908_7d5c_f1b0_2fec_b556_2e02;

        #200;
        key = 128'hdcda_4650_573d_0f94_f934_add9_5ae7_3b2d;
        state = 128'hbf29_b616_d5c2_5b64_315b_5d70_8d91_ffa2;

        #200;
        key = 128'h926d_f192_3313_1a34_4cd5_715c_0695_e66f;
        state = 128'hd054_1c91_c129_8ae0_1a28_5431_1567_f4e9;

        #200;
        key = 128'hebe8_5fa4_e8a4_d2b3_e606_c03a_4259_9127;
        state = 128'h02b2_b550_e357_9533_50a3_0121_3f5b_2b5b;

        #200;
        key = 128'hbe20_928f_5faf_3bb0_2701_da8d_9059_5e4b;
        state = 128'he3a2_3f88_9b36_f7cf_bea8_b918_0442_517c;

        #200;
        key = 128'h2097_60ab_b1fc_13e2_bed0_204b_b530_bb79;
        state = 128'h1114_6cd0_c2cf_a485_cb35_f773_bd24_9381;

        #200;
        key = 128'h65d2_df99_0f83_073b_c42c_da84_1733_b5a3;
        state = 128'he4ce_64d7_5fac_29a8_2387_ce6d_1ac2_8445;

        #200;
        key = 128'h44fc_962f_8be6_4084_43b6_77ee_5b06_d223;
        state = 128'hb308_2383_e484_2605_76ca_7b20_7d85_05c6;

        #200;
        key = 128'h7787_28c4_34fc_c290_1183_5f0d_4c33_abd2;
        state = 128'h373f_df37_0a79_2e67_b6dd_ca54_ad47_6e82;

        #200;
        key = 128'hec39_db42_7c08_5b68_1e1e_cf03_817f_327d;
        state = 128'h348a_33b1_3235_e18b_28a2_7ab6_35ea_5236;

        #200;
        key = 128'he96c_aa65_6bad_03b5_9079_d233_40e7_52ad;
        state = 128'h59d8_3e02_7030_d064_79c4_f143_6e21_53c8;

        #200;
        key = 128'h0454_cba1_444e_80c4_f0a4_6b06_4f80_a1f5;
        state = 128'he432_6f14_4ac1_1281_f5e8_f593_7069_4c47;

        #200;
        key = 128'h0033_f51a_765a_4668_9568_f821_1d62_22c1;
        state = 128'h8ef9_ddb1_7ba9_64f8_27e0_ab46_967f_6f56;

        #200;
        key = 128'hbfcd_a779_56c5_c981_5420_567a_94e5_a9c5;
        state = 128'hfe17_f215_332c_1afc_82f8_a5cf_4f77_a6be;

        #200;
        key = 128'h7940_0986_d767_5792_f0bf_8cd4_12a1_087f;
        state = 128'ha843_a306_9588_7f37_db35_1e9d_5f7b_39cc;

        #200;
        key = 128'h9558_7b3a_0c7e_a560_80c9_25e8_1ec8_90a9;
        state = 128'h400a_b5b7_9928_1a88_45a9_4a9b_d2fc_a239;

        #200;
        key = 128'hc33a_5350_4280_87c8_2ff1_da49_37b3_d2b8;
        state = 128'h41ee_da44_cf9e_b201_49d6_6628_91a4_89de;

        #200;
        key = 128'h3fb4_d9b5_8997_d824_d697_fc2e_d557_2586;
        state = 128'h97ec_cda8_bd45_15f6_603f_8d98_ea84_6ce0;

        #200;
        key = 128'h9334_ef27_24e1_5acb_c6d8_9c70_ae33_2edd;
        state = 128'ha718_cbb7_6de8_7aba_881f_c181_916d_5911;

        #200;
        key = 128'hfbea_19b0_b62a_83b2_70f9_7f76_3a7b_cec2;
        state = 128'h6c7b_6a7b_53f5_32fb_21d8_7752_9dc4_e13c;

        #200;
        key = 128'h54aa_b404_134d_4621_b780_c650_708e_4ac6;
        state = 128'hecd0_4961_5c65_3c91_788b_0d68_fbe1_6df4;

        #200;
        key = 128'hee6f_a7d7_e615_fc39_fcdf_218e_fde4_e02f;
        state = 128'h9baf_7a54_542e_28fd_8181_f72c_b313_cc27;

        #200;
        key = 128'h57af_f8a8_a7bc_3d76_2ae6_6c22_8149_7052;
        state = 128'h7363_007f_4638_17d4_e704_9362_b9fd_80c6;

        #200;
        key = 128'h41ed_46d5_4412_4f16_1baf_4f25_fd9b_4405;
        state = 128'h1987_8043_c9e7_9d85_f5eb_ed61_0a8c_facf;

        #200;
        key = 128'h1238_7ac5_99fb_3182_2a8a_8efd_b405_8e94;
        state = 128'h7656_2f5f_b0b4_01f6_5411_658a_d79a_622a;

        #200;
        key = 128'h56e1_0813_b1be_0e07_9895_3725_d73b_709e;
        state = 128'h2a8b_c1b1_9119_e562_25fe_2e7e_6e45_f9a6;

        #200;
        key = 128'h00ac_e6b4_2aac_5f01_6d04_89e5_5f03_4773;
        state = 128'he4df_4136_6181_d3c3_3ed5_4ca8_64af_1566;

        #200;
        key = 128'hef8b_b03a_ede8_fe80_2d3c_bda8_e995_0001;
        state = 128'ha7c3_9e96_6078_58c6_ad2b_1724_489f_42aa;

        #200;
        key = 128'h2e61_9261_b2d6_011c_69fb_f937_0abd_6e2b;
        state = 128'h550b_f238_72e2_513d_785f_27a5_3351_3c75;

        #200;
        key = 128'h9258_8e59_3b2c_dfeb_feac_359e_a1ec_75f6;
        state = 128'hc6d1_cda9_0a93_5cc5_2628_3103_1295_7b4b;

        #200;
        key = 128'h8a48_e3f4_fa09_6d44_88c4_edaa_5614_72ec;
        state = 128'h5896_f302_982d_e835_dbe5_af3c_d5c0_4c83;

        #200;
        key = 128'hccce_a598_6745_c28e_67f5_ee82_9ba5_6656;
        state = 128'h0581_2d43_cdb7_9d1a_8b9a_3cd6_8a8f_1bb7;

        #200;
        key = 128'hc44d_e529_4605_766d_1f87_7fbe_96ff_0d0c;
        state = 128'ha804_70d4_a810_5548_6361_eeaa_88d4_0e93;

        #200;
        key = 128'h678a_48be_f3d7_7130_dcac_7725_aaae_401c;
        state = 128'hfd25_e465_66af_7ca9_85ea_cead_f549_77fc;

        #200;
        key = 128'h2277_bbe8_e5f8_72be_e8d0_84dc_b67b_e9c3;
        state = 128'h9d4a_ef16_c371_3eef_09cc_e4bb_47f2_a60a;

        #200;
        key = 128'h19b5_b985_4663_1fa3_5b57_a1c8_4fe4_dde0;
        state = 128'h9aa0_66a0_f755_88c8_169a_0166_7f44_adf0;

        #200;
        key = 128'hf139_ca26_409f_4d8b_c343_10e1_e928_9f09;
        state = 128'he17c_16ad_f5d8_259c_177e_5510_c910_81af;

        #200;
        key = 128'h93f6_2d83_64d0_5657_9a7e_065b_2f1d_aa45;
        state = 128'hfe57_2087_7ac5_e608_3ae8_24c9_e893_c713;

        #200;
        key = 128'ha9aa_ab4a_197f_b032_d88f_7e4d_305c_15cb;
        state = 128'hd984_fad8_2ce9_e983_4d99_8a6f_c3ba_cd50;

        #200;
        key = 128'h9bbf_ddcd_c0e4_6eec_3f18_1bbd_4ad1_999e;
        state = 128'h34a0_a9dc_38f7_3b59_4136_8a23_f137_a50e;

        #200;
        key = 128'h34d6_38f7_5779_ee26_57b9_5182_6b3a_ea2d;
        state = 128'h2e2e_4878_27de_b499_cce7_1e94_1320_a6d8;

        #200;
        key = 128'h8e1a_661c_8681_f76d_5012_4840_70f5_e533;
        state = 128'h60fd_1c3e_a3dd_aa29_37c6_9ccc_7ae4_1e58;

        #200;
        key = 128'heda7_aaa4_962f_33de_8feb_b484_e682_dc9e;
        state = 128'h61ab_1a22_993f_1da6_02d0_6ab5_e359_6517;

        #200;
        key = 128'hbc45_9a3a_e59e_b2bf_03e0_0d4d_3bfc_b107;
        state = 128'ha581_64c6_4541_a426_9591_345a_e7dd_8e32;

        #200;
        key = 128'h65ef_fc15_e41e_39e2_40e4_332f_bb3b_b81d;
        state = 128'h5bcc_a0dc_accc_468b_bed2_35db_e4cc_8084;

        #200;
        key = 128'h9f3c_b70b_d81c_bc35_f255_c5f4_f0e4_6754;
        state = 128'h2284_b551_df16_d65f_80ef_cc39_04e3_6aa4;

        #200;
        key = 128'h21b4_7552_b0ca_ea69_9e39_7da6_ec12_d368;
        state = 128'h98f4_9e96_168b_f74d_7958_e349_2b11_7631;

        #200;
        key = 128'heef2_5a8e_d3ee_c6c4_31a3_7974_e485_b0da;
        state = 128'hc2ce_e1f7_aa6e_763d_70d8_4099_316c_bd75;

        #200;
        key = 128'he47e_f6a0_fefe_25fb_0e2a_e153_2171_1312;
        state = 128'h82d9_ac97_33c3_0c6c_72aa_d9c7_4e7f_23ff;

        #200;
        key = 128'hcaa2_4fd4_d2ac_fa69_b04d_de5d_17a4_75ae;
        state = 128'h9c88_6edd_c87f_21e9_22cb_99ae_c9a4_9f09;

        #200;
        key = 128'h9617_dd80_cb75_b364_d2f0_1548_203f_3c9d;
        state = 128'h0a59_3d49_2b3d_5764_08bc_2d81_5790_fa84;

        #200;
        key = 128'h343e_f6fd_1fa2_8e5f_0ea7_712a_30b6_7b3f;
        state = 128'hf135_12b9_369e_a3be_2238_a9d3_5f8d_7dca;

        #200;
        key = 128'h79f0_4a90_fd27_e79f_ced7_78bd_f2ab_fe03;
        state = 128'h877b_dc92_50c0_d129_9645_8ca3_d08a_29d2;

        #200;
        key = 128'h173d_4542_5864_1bbc_ec8b_2720_7643_2113;
        state = 128'h2368_52ab_656f_8d34_6e05_5f09_b6ad_4e13;

        #200;
        key = 128'hcc90_64b8_ba8d_dfd5_e921_82a8_5929_8a14;
        state = 128'h94f0_523d_3705_166d_fb34_14d7_ffba_5454;

        #200;
        key = 128'hadfa_e492_ce6d_0339_c7b5_3293_a665_5293;
        state = 128'hc467_d77f_5f6b_ccbf_d9e2_7fdd_f0b5_54c0;

        #200;
        key = 128'h2494_68f9_7282_91e2_5b2a_c92d_ba60_a2e5;
        state = 128'hbbd6_2283_a602_2ffd_48ae_9739_fd85_cdc8;

        #200;
        key = 128'h6804_1f51_dbc5_bd81_620a_0955_1871_dcdb;
        state = 128'h72ee_51c8_5a77_baa5_249a_8312_69aa_0b2c;

        #200;
        key = 128'h08ca_0b4d_c75d_98ca_e5a2_5dcf_5c83_2a63;
        state = 128'h1a4f_23d9_df4f_9e62_56c3_3b44_f13d_e5c6;

        #200;
        key = 128'he4e5_68f0_581f_5b24_44c2_9669_6975_508f;
        state = 128'hcd9b_26e7_433b_e8bd_b65d_b4b8_e017_379c;

        #200;
        key = 128'h2333_9c6a_fe0a_9ce4_bc1e_b3b0_4e85_6f4d;
        state = 128'h0d1e_ff41_ec30_7d26_b274_774a_cab1_0470;

        #200;
        key = 128'he9a4_8bc1_113a_1498_4bce_2955_3cfb_f1e0;
        state = 128'h7652_bd38_afee_e4e6_3cb7_c9ec_5238_ec7c;

        #200;
        key = 128'h0acc_126e_e4fc_1acc_6daf_1378_9d3a_b582;
        state = 128'h3def_bca5_635d_70ad_ac61_78c3_d9f2_a2dd;

        #200;
        key = 128'h077d_671d_29c3_34ef_5856_02cd_ace7_4749;
        state = 128'hf645_257d_4fa7_0e6d_0999_5342_65a4_93d6;

        #200;
        key = 128'hea1b_b564_d973_7a2a_2ff8_b99b_c4fb_c865;
        state = 128'hc1ae_1992_85ed_96ae_2a46_d05f_da59_b955;

        #200;
        key = 128'h64d9_5a90_8a69_f449_1bdf_a947_4674_2799;
        state = 128'h0930_99e4_51ac_569b_3243_1a62_2fb9_6341;

        #200;
        key = 128'h0d76_9f17_313c_e74e_1e71_018f_c228_076d;
        state = 128'hc343_7748_41ac_c605_940b_1fa7_bc01_b1a3;

        #200;
        key = 128'h5c1c_2610_09b1_48ea_fed2_5ef2_856c_8b4c;
        state = 128'h3a3b_964c_1e1c_e9e3_d36b_d761_4b7a_560d;

        #200;
        key = 128'h12f7_b9e8_2783_c73c_1f8e_2d35_9e9f_8731;
        state = 128'h7bc4_0b83_41c1_50ac_98d5_4cfd_f4f0_4e7b;

        #200;
        key = 128'h4a25_37a6_a0aa_69ed_a661_b963_4ef8_fc9e;
        state = 128'hc2b2_9141_5b34_5c9b_f149_ba94_751d_1753;

        #200;
        key = 128'h298c_0198_2f4f_f85a_050e_87e9_cdf2_21bb;
        state = 128'hb875_8669_1bd7_8a83_b0c3_4c63_726e_d314;

        #200;
        key = 128'h5fd6_c611_7331_fbdc_ab9f_5bd2_deb1_530d;
        state = 128'hf79b_5627_0146_8211_e8ad_2aef_08d9_efef;

        #200;
        key = 128'hfb84_7dde_bf1c_28e1_d71a_3755_25d0_da67;
        state = 128'h63d8_378c_7ede_c79f_8799_bb89_ce37_1a0e;

        #200;
        key = 128'hc34c_d78b_2b3e_b940_9485_0d7e_4047_bacc;
        state = 128'h7d53_9537_9bc5_bf41_881f_8dc5_5dac_a409;

        #200;
        key = 128'h8f50_5a8c_67ac_4955_c590_8d1b_71dd_33ab;
        state = 128'hcdeb_d04c_459c_026f_26b3_b9e3_54a4_1f32;

        #200;
        key = 128'h74a0_b4a6_eeee_bf21_e8e7_5125_22c5_2d67;
        state = 128'h5dc2_aebe_4ea0_74dc_9304_ea00_5f13_dd0f;

        #200;
        key = 128'he04f_c535_7bb8_4b7c_0a4f_b59f_2d3a_4146;
        state = 128'h835f_6998_965e_29f2_d40d_c7b0_84e5_a3cd;

        #200;
        key = 128'h5751_eabe_d8de_536f_6e1f_a047_49ce_4dbf;
        state = 128'h64ed_4754_dd5c_248a_85d5_da71_cef9_769c;

        #200;
        key = 128'h54bd_9cc5_80f9_133a_f203_9c28_4782_26ed;
        state = 128'hef52_3628_3215_543b_1a26_c0c3_d609_fcf9;

        #200;
        key = 128'h5c82_4015_1ea9_99a8_9ead_b20f_9729_6842;
        state = 128'h3335_df51_da54_fb81_565d_391d_06b6_2e48;

        #200;
        key = 128'h88e0_9c04_8e46_ecfd_6b0d_e5b6_010c_8a2d;
        state = 128'hf7b7_156d_6f6b_1017_8503_2227_2921_f359;

        #200;
        key = 128'hdac9_a413_7417_6b6f_1db3_17bf_c509_5b12;
        state = 128'h1771_a6ae_5124_5d85_2716_fa3f_012d_3f9d;

        #200;
        key = 128'h6e9e_0790_0c51_08d8_08d5_be4a_3d8a_eb59;
        state = 128'h37da_906d_31f0_2658_afd5_2503_0f38_f912;

        #200;
        key = 128'h0bc8_d25f_f89a_4569_8010_b8f7_cb1f_696f;
        state = 128'h1928_5ebd_c237_9675_c305_24ac_857e_3b8b;

        #200;
        key = 128'haf0c_1115_0d1d_9a18_e390_4538_27e1_b52a;
        state = 128'h8175_0c33_9f36_3f2b_10cb_82d3_3ab0_df40;

        #200;
        key = 128'ha5d0_9542_f97a_3754_a35c_fda0_6128_8406;
        state = 128'h6d5e_0ed0_3faa_0adf_7b62_dfa6_3759_7edb;

        #200;
        key = 128'h973f_0667_ac2e_e3e4_95c2_87d7_a1fb_7d58;
        state = 128'hf752_c23d_5d43_f293_d25c_2242_04d2_b028;

        #200;
        key = 128'h2fcd_44ba_a71a_b149_115d_d325_36ff_7d5d;
        state = 128'ha077_7425_3efa_ada9_6534_899d_8d7e_5cf5;

        #200;
        key = 128'h8aca_a5fa_3205_d4a3_cc1c_b003_3571_2401;
        state = 128'h2067_032e_b5d7_ffda_2270_ea5d_4d8b_5232;

        #200;
        key = 128'h541d_4c10_18e2_fd15_b0ad_b6eb_3a94_5e70;
        state = 128'h4297_45e2_3704_bb99_c37c_8179_a31e_3433;

        #200;
        key = 128'h8be5_7791_adb9_09a9_1b05_75d7_17b9_0c23;
        state = 128'h5abe_3570_a460_07bf_60f9_4a2e_169b_6ba2;

        #200;
        key = 128'h06aa_6f39_96ba_b45e_6b48_2d08_20bd_d7d4;
        state = 128'hf516_9545_444b_bae5_6087_0445_5991_2b00;

        #200;
        key = 128'h0e66_be8d_0038_8230_1a39_0970_eef7_6288;
        state = 128'h95f8_5e09_9dea_6c8d_4686_80e3_e931_fd50;

        #200;
        key = 128'he5b1_426a_04e0_706f_8189_16b8_36d4_d6f1;
        state = 128'h5568_fef5_ca78_f020_0eb1_20dd_4d69_a3b6;

        #200;
        key = 128'hdd9b_08c9_1376_6368_d4ad_5953_a9c2_6be5;
        state = 128'h3716_57b4_9c5b_6aa8_31b8_dfcc_4a82_59e4;

        #200;
        key = 128'hd59c_356c_b5cd_0f14_0481_c648_92af_2788;
        state = 128'h4a96_307b_d1b0_40b5_a9a5_87c8_42e5_271c;

        #200;
        key = 128'h1e9a_8546_20cc_23db_55ca_193c_c59a_256a;
        state = 128'h2c96_f168_125d_b8c7_93c3_8ec2_885c_5ba1;

        #200;
        key = 128'he7b8_a080_1f7e_d137_7e89_8227_b511_012d;
        state = 128'h01e4_fe9c_61a5_ce3a_d130_5647_bc87_ddcf;

        #200;
        key = 128'he56c_1f36_247e_67f2_6af2_c99b_cb28_8473;
        state = 128'h34cd_a202_b3d3_bbb0_ff93_e273_900a_605f;

        #200;
        key = 128'h8e73_e90b_ae14_bfb4_22bb_cd32_d2d4_27bc;
        state = 128'h399a_d5f9_d2fe_a9cf_aa9c_215e_774a_3474;

        #200;
        key = 128'h5787_0320_0ebb_1b78_fc27_e4ab_81a6_2d5a;
        state = 128'hd1cb_bca3_87f8_083a_d620_cc05_6923_e752;

        #200;
        key = 128'h1695_4303_99c4_41f7_8e1c_a511_aa72_291d;
        state = 128'hee83_bfee_ca04_7882_1e6c_b2ef_8528_6269;

        #200;
        key = 128'h0fa0_18c3_6d9a_ea7e_eeb9_ad1c_5f5e_5c81;
        state = 128'h29ae_0465_1247_8431_13dc_225d_e1fa_7fd7;

        #200;
        key = 128'hd093_16a6_6763_2bab_dc40_d3ad_dc09_3654;
        state = 128'ha16b_48c9_91bf_f746_1216_1a4b_6941_a1d9;

        #200;
        key = 128'hd061_c471_7dca_5937_8937_ff5e_fb56_cd70;
        state = 128'hc5f4_40fd_fb72_095a_35d4_4325_455e_8fa3;

        #200;
        key = 128'h700b_4c78_6ff4_f61a_110d_d53a_012e_3b8b;
        state = 128'hdc54_b8c5_458c_10f4_83fa_6d22_a08b_fc79;

        #200;
        key = 128'h8ef9_e7f8_20d7_9c2d_db17_08af_af49_97a4;
        state = 128'h264d_bc7c_cc6b_f100_6413_5668_da8b_c133;

        #200;
        key = 128'h6581_dd99_ee8b_2e90_6fd8_597a_36a7_ab61;
        state = 128'h545e_e450_4a9b_d050_7cde_b552_ad65_398f;

        #200;
        key = 128'h399b_6594_a63e_62fc_5eca_60fc_e1a6_6c0e;
        state = 128'h651d_02c7_4cbb_a245_5e95_0ef2_6cde_efff;

        #200;
        key = 128'h0f25_3ed3_b366_7645_a6b6_1652_b96a_3eea;
        state = 128'h4e12_5708_09b1_f91c_93cc_3967_2e69_3e02;

        #200;
        key = 128'hd784_9cc9_4c5f_9cf9_4976_2f55_d3ef_9968;
        state = 128'hd290_f2b8_7329_0092_da53_58ef_d810_1808;

        #200;
        key = 128'h563b_9bb5_d8ed_d963_29b7_64ce_9bac_5e54;
        state = 128'hee0e_63ae_d228_30cd_8dcb_d2ce_e1a4_c6cd;

        #200;
        key = 128'h2cd2_4654_042f_7348_3651_5712_4cd6_020a;
        state = 128'h9592_1d38_c9a9_e110_5ac9_fc5f_22a0_c8a6;

        #200;
        key = 128'h2a40_96c9_d294_647b_2747_e6e8_93fd_9a81;
        state = 128'hcb06_15fd_28a7_25e9_883d_bdb1_b42a_4c11;

        #200;
        key = 128'h2097_39ea_1b7f_ead7_bac8_0813_6c4e_57a2;
        state = 128'hf0b7_4af9_3880_adbc_28f0_61d4_8da6_5dc8;

        #200;
        key = 128'h737f_2d67_1d5a_8b29_609c_362b_c11a_8a49;
        state = 128'h3a7f_392a_0473_477b_7f5c_54a0_c2da_64a3;

        #200;
        key = 128'h37c9_d600_5612_45ab_1935_c99a_9ba3_e5f3;
        state = 128'ha1cf_bf62_5707_4cc7_dec4_5dba_939a_03f9;

        #200;
        key = 128'h4403_f808_d3f7_20c8_af82_1552_2304_7d7c;
        state = 128'hcc00_841f_15a5_ff26_e593_45aa_8008_f5d6;

        #200;
        key = 128'h37c6_91a0_252b_8f49_aae2_e55a_9881_b75b;
        state = 128'hd5ae_1389_34d2_424a_6829_21b4_ee2e_8ef7;

        #200;
        key = 128'h226c_1c7d_c1d3_16fa_cc8f_62de_94ab_3798;
        state = 128'hd557_5ef0_b30f_961e_e089_47da_a3d2_e558;

        #200;
        key = 128'h5777_ec65_1631_9a8b_8989_4543_970d_eaff;
        state = 128'h4696_1c7c_ea55_b302_a4f2_f1aa_d8e2_c88b;

        #200;
        key = 128'h0c39_ed4b_2081_b374_3355_ebcf_518c_c9f2;
        state = 128'hb444_30f5_4825_d635_26c4_d1d6_85bc_e652;

        #200;
        key = 128'he889_cf60_c748_276d_9ca1_842f_1583_fdf7;
        state = 128'h0f49_f2b8_b55f_f726_e171_d06d_b03a_ee30;

        #200;
        key = 128'hd9ab_6d31_937f_cb7a_e136_bf85_49eb_d0fe;
        state = 128'h8ffe_5c25_9060_c843_ccd3_2884_c188_73ba;

        #200;
        key = 128'h74b2_f003_4f05_26ee_8966_a059_9455_5fc2;
        state = 128'ha25d_44ed_78c9_eeaf_c2ff_f8b6_db13_872b;

        #200;
        key = 128'hdb7b_b99b_7abd_a58b_20f5_a13f_7f5d_11ec;
        state = 128'hce53_6b80_1ceb_96f3_9c74_999e_5b21_7d01;

        #200;
        key = 128'ha4f1_0802_6218_3644_55d2_97f6_25fa_6449;
        state = 128'h0982_d135_182a_5fba_3ac9_b47d_a0bc_ba9d;

        #200;
        key = 128'hdff0_a401_225b_5a95_5ef8_e999_eeb5_c6cd;
        state = 128'h3107_91e3_3d36_7c22_b8ab_851f_2b65_5cf9;

        #200;
        key = 128'hcef4_d16b_f133_9b7d_7eed_320f_459c_509e;
        state = 128'h1af4_f586_24f2_0038_300a_02f8_7b4b_696b;

        #200;
        key = 128'h39b8_f4f7_f743_1cf6_e994_47d1_b259_f8d6;
        state = 128'had33_c592_8a05_f7ae_6e41_dbdb_9b61_1732;

        #200;
        key = 128'h370a_1dda_c7f3_1eb1_6800_35a5_d22f_8c65;
        state = 128'h442f_5041_55e2_a01b_4b82_e963_2f15_14bd;

        #200;
        key = 128'h7b14_a1a5_d923_14dc_9dba_658b_b3b1_d340;
        state = 128'ha4ec_f2e0_39dd_8f29_9eaf_a2bc_e97a_de33;

        #200;
        key = 128'h01e7_b130_feb5_bbad_0421_bdc1_8e2c_0270;
        state = 128'h850e_12a0_dfda_c0bd_0caf_fe90_e0b6_c52c;

        #200;
        key = 128'h6c6c_8efb_3237_b299_4cc7_4fb7_5bbc_b04b;
        state = 128'h83b4_45cb_65bd_8a90_da88_2a21_6366_43d2;

        #200;
        key = 128'hf812_9671_13c8_f7cf_570a_f811_aacd_2107;
        state = 128'hdb40_c4b1_69c0_631b_4e85_fdce_1e79_5e50;

        #200;
        key = 128'ha48e_0b52_88db_a3ae_de4e_8243_6c23_fb4f;
        state = 128'h29db_3715_b844_6fac_8a1a_c24d_79f9_6391;

        #200;
        key = 128'h2608_6086_4439_7c75_7994_0df0_295f_d1d0;
        state = 128'hbcdd_1f0f_e0d6_721c_a2e5_12da_1bec_c7a6;

        #200;
        key = 128'h5813_a5b4_b7fd_7e52_030c_6c80_9d08_b7e8;
        state = 128'h8918_9c40_5832_cd56_464d_e7e6_66b3_6c86;

        #200;
        key = 128'h906b_02fd_e6ca_e99e_5f80_5191_76c6_c963;
        state = 128'h7c8d_7bf2_2b8e_587e_5a08_68c8_d89b_3221;

        #200;
        key = 128'h77c9_8969_3df7_fcd5_1024_f6a5_0e6e_f11a;
        state = 128'h00a7_85e6_636e_69bb_3ae4_e9af_c50f_68be;

        #200;
        key = 128'he71b_cab9_8649_dca1_f322_6dab_2f2d_85f1;
        state = 128'hcbc1_89ab_f4bc_6092_11b3_faa5_683f_f274;

        #200;
        key = 128'h799f_ac9b_e9c6_a9f4_1e9d_fe24_5b12_e8d2;
        state = 128'h2750_ef91_a653_4310_efa0_0688_67e4_38f1;

        #200;
        key = 128'h45e9_5e45_03ec_43c7_fae1_95bd_2dd6_43af;
        state = 128'h8e89_34fd_4801_a715_19e0_fab7_233b_6096;

        #200;
        key = 128'h8392_dbd6_b1b4_51ea_cff9_483c_09d8_9eb4;
        state = 128'h9cd4_7c74_e6fa_e6d4_d133_1a79_6483_2fc3;

        #200;
        key = 128'h496c_6d31_86c0_6856_15fa_fb0b_ad73_fe30;
        state = 128'h52be_f492_d8b7_7006_8ed6_83ca_cec3_3011;

        #200;
        key = 128'h23fe_e9c1_cfb2_7a2f_c720_09c1_e6f9_85ee;
        state = 128'h868b_1e3b_4282_d872_92a8_2c57_5d65_213d;

        #200;
        key = 128'h0217_3aeb_ffa5_f059_d1fc_d623_c6e7_fdda;
        state = 128'hc03a_6357_e47c_ae5d_507b_c815_2c19_01a1;

        #200;
        key = 128'hee7e_3cc9_316d_bd2f_4c15_382d_d923_3a58;
        state = 128'h71a7_a3bd_886d_0204_180f_0ff1_a5c0_f699;

        #200;
        key = 128'h855e_5ab1_ff21_235a_288c_31f4_cd1d_49b7;
        state = 128'hb520_3cc1_2fbb_67b2_bb38_6266_757c_53b3;

        #200;
        key = 128'hcbf4_6812_14c2_17e4_6c8b_ca19_985c_c6a2;
        state = 128'ha023_e2d5_d8dc_fbdf_d232_e791_e84a_c328;

        #200;
        key = 128'hd514_21b1_a8bb_b288_9635_b053_6dac_11e9;
        state = 128'h7804_aad1_5412_6a79_b41e_9f48_895c_345d;

        #200;
        key = 128'h75bf_befc_4a08_5949_2e91_44aa_e8c2_cbe1;
        state = 128'h6dce_0d69_dd98_8011_cd9a_c092_e0b0_29bc;

        #200;
        key = 128'hf9e2_436a_2be2_b4a0_abed_ca79_5c59_9902;
        state = 128'hedb0_5b0f_4123_7660_2e34_8ac0_8235_8b51;

        #200;
        key = 128'h5722_bc09_12e2_ca57_740a_8e1e_2988_0831;
        state = 128'hce14_81ae_5202_3f83_b5f4_1437_8fc4_645f;

        #200;
        key = 128'hc5d7_dd1d_66ca_e455_830f_6f94_2094_eb61;
        state = 128'hd1d7_e362_98e8_cf52_2bd0_d1b1_6d96_1f27;

        #200;
        key = 128'hb525_dde8_b0ba_b7c3_0703_f6ac_9d28_72ff;
        state = 128'h0b3e_6929_6e64_e898_3e70_c44d_6bad_39e1;

        #200;
        key = 128'hdf7d_9627_2336_7399_93aa_72d8_c9b1_e69a;
        state = 128'h0a45_aec9_4f49_6d82_6ca1_d916_07eb_50dc;

        #200;
        key = 128'hc4a5_0cae_7a19_413c_9001_fef8_2e90_486b;
        state = 128'h5ccc_e2e5_5019_47ba_088d_7453_64ec_3fde;

        #200;
        key = 128'habce_5cb6_9d8b_b87d_c4d6_bd52_4f0b_8de8;
        state = 128'h5236_7a7b_f54b_27b2_c43c_2298_cea3_c9b3;

        #200;
        key = 128'h5d61_7fb0_ad08_dd11_123c_0adb_e4ed_9fc9;
        state = 128'hc0f3_33d1_92ea_658b_5ae9_ad20_ce2a_8d63;

        #200;
        key = 128'hb545_a196_38df_02a7_30d6_33bc_ecdb_336d;
        state = 128'hc8c3_a12b_e698_5ea2_ce8a_8886_ad2b_39a7;

        #200;
        key = 128'hcd66_0a01_7603_c363_bf43_b556_3a69_bedf;
        state = 128'h9fe1_7e91_c628_7dc8_8899_0bbc_f6a4_e83e;

        #200;
        key = 128'hdecc_8a72_7199_98a6_fc43_7ec6_837a_3f16;
        state = 128'h3f28_cc77_f4be_0f1e_a99c_b27a_748c_a89e;

        #200;
        key = 128'hd1d2_a67a_299b_7d01_245d_a79e_6fe0_9441;
        state = 128'hac0b_8f1b_1b36_52fb_64a6_959c_12ce_f30b;

        #200;
        key = 128'h8a37_3860_46c1_56f1_c363_1f00_d21f_5e96;
        state = 128'hf7ff_a792_160f_52a2_2d52_96d7_097c_dc6e;

        #200;
        key = 128'ha77c_1122_637a_448d_98a8_dafa_6fc7_7bcf;
        state = 128'he96b_cb34_195c_4b69_c50d_de3e_32e0_1b20;

        #200;
        key = 128'hbb33_5d42_0d49_fa59_01ec_1bd0_d68c_f1d5;
        state = 128'h5ac0_3c51_af8f_81b0_6637_be35_34d4_09f7;

        #200;
        key = 128'h9a61_5920_0764_5373_2c88_878f_f892_e231;
        state = 128'h15d9_51f4_c2d4_fb6c_eb83_f5f4_bcef_f896;

        #200;
        key = 128'hcff8_bffa_6cd3_d06e_83f6_4d56_ce7d_c0fc;
        state = 128'h865a_4119_b18f_59b0_bdf0_7300_36c9_afb0;

        #200;
        key = 128'h89ea_4baa_047c_7143_d4f5_b9ae_f8d6_72ba;
        state = 128'hbdbb_ab81_c7d8_d869_f229_6df7_6326_3167;

        #200;
        key = 128'hd7d5_aa4c_ac6a_4d39_c768_72b7_e8a8_4db6;
        state = 128'hf068_9ed1_68d5_6a1f_77c9_3657_744f_7502;

        #200;
        key = 128'h8f82_4b4a_d374_dfef_2bd6_7a74_91f0_a8e5;
        state = 128'h472c_1289_00dd_180a_13f5_f3ad_2a89_c00d;

        #200;
        key = 128'hab7e_a3ba_68e8_439b_8820_8a00_8645_1c3c;
        state = 128'hd0da_8d1f_4085_b976_a755_2721_0db8_5e86;

        #200;
        key = 128'he7ba_4e38_d2e4_6e57_d4f6_d318_a556_38bd;
        state = 128'h034b_a5d2_1833_100f_3f5b_8542_0ce5_ff60;

        #200;
        key = 128'h7fc4_bf41_66be_6b04_7030_ce6c_205c_b7da;
        state = 128'h868d_95f4_70a9_71ce_edbb_141e_97c9_643c;

        #200;
        key = 128'h5fef_4bb2_642f_d310_8916_89fc_6f05_ab7b;
        state = 128'hc68d_c75e_1b8e_2bb5_399c_de80_da76_f93c;

        #200;
        key = 128'heae9_16c9_e2b3_c22b_a857_3df6_5cdb_0ee4;
        state = 128'h1713_95ca_e073_f3af_fdfb_67b0_c432_d352;

        #200;
        key = 128'h05a0_015c_d02e_df5d_0cfd_2f9c_1fd9_c9bf;
        state = 128'h246c_bbe3_a42f_3e65_11c9_0ee8_fdd3_3d84;

        #200;
        key = 128'hedd9_6e3f_876a_b1d4_e400_fb4f_525a_45fb;
        state = 128'h4c1a_6e62_460f_e57d_78fa_6e71_514a_91ab;

        #200;
        key = 128'h2073_ce91_620c_8ec2_decc_0b8d_f73d_79f6;
        state = 128'h7cde_b21f_2b71_6a9b_d3ed_a7ec_8c2a_314b;

        #200;
        key = 128'hf30d_24f7_9f27_da04_df34_072f_9293_35ad;
        state = 128'hfde5_c5bd_c0bf_9975_887e_cd24_44c4_57a3;

        #200;
        key = 128'hbc60_25d7_38fb_cd14_dcf3_4964_c49d_aa8e;
        state = 128'h5f4f_487a_51af_35e2_8f94_26af_d646_da19;

        #200;
        key = 128'hd3ed_f4e6_e5d4_2eb5_58aa_db93_6a2a_0628;
        state = 128'h5559_8e90_4e90_a336_f680_ecb2_4826_e452;

        #200;
        key = 128'ha1ae_ce6a_2d0e_2cc9_4ba7_2af4_15a9_7320;
        state = 128'hb5d1_5095_acc8_db77_3110_5cb2_b629_254d;

        #200;
        key = 128'hd304_d988_f369_69e8_f5a7_1f86_e1ee_28df;
        state = 128'h184b_22b6_d9ae_c92c_4111_011d_ea73_27db;

        #200;
        key = 128'hcf60_7ce2_a8cc_fa27_33fa_eeb9_6cbd_fabb;
        state = 128'hee80_b9c6_386c_887c_544b_32d4_aa0d_9c45;

        #200;
        key = 128'h2b2a_80d7_66fc_8ded_dd16_ceea_93ab_8123;
        state = 128'h9496_f9f3_e091_9510_5a22_30ef_5020_d9d5;

        #200;
        key = 128'h305c_e683_1fd1_4ed4_6785_fa2e_02e6_e137;
        state = 128'h05c1_6cc9_dd41_e86e_e510_fde8_21f3_7531;

        #200;
        key = 128'h6674_1d5d_4335_5e5f_bfdc_7510_c9c3_134f;
        state = 128'he6ee_d4e4_464a_2e81_1785_c215_b646_3495;

        #200;
        key = 128'h8fb4_e3af_f5b2_545c_e289_5bd6_e923_5176;
        state = 128'h182d_1334_ee63_e954_d388_c762_93b6_80b3;

        #200;
        key = 128'h5481_9a60_f3de_1e6f_47be_6a46_7d7a_dc39;
        state = 128'h70a3_f25f_4268_d09e_65b2_72e8_91f4_67c9;

        #200;
        key = 128'hde30_34b9_1d4d_d8f8_b606_59a1_90d4_bc4e;
        state = 128'hde5f_d106_54a0_a77b_c258_e275_552a_7914;

        #200;
        key = 128'h3856_848d_235d_adef_0818_93d5_3bd4_f8d9;
        state = 128'h0e65_3734_87bb_5aa1_ff63_2293_a407_6b28;

        #200;
        key = 128'hdad2_c233_ed10_9876_9a3c_91cd_26f5_4ffc;
        state = 128'h4509_51a2_1af6_7628_5b7a_3c55_5221_8e3f;

        #200;
        key = 128'h0b83_59ea_92c4_2175_f013_504f_20be_f68c;
        state = 128'h3e09_d04b_fc53_8806_b757_2e89_7ae1_ed25;

        #200;
        key = 128'h2875_4c26_ed3c_602c_7d83_acaf_31a8_c6c0;
        state = 128'h9320_b56e_ef18_dde5_e664_6a55_429c_4b89;

        #200;
        key = 128'h3e89_54c2_ddac_e37b_ea72_19d8_7d82_ece3;
        state = 128'he6a2_4239_1a94_01f0_f585_55f9_f7fc_0ef2;

        #200;
        key = 128'h312d_17c9_a7bc_ed69_f125_dd99_3173_3745;
        state = 128'hf263_1806_b0ef_ea44_d2e0_8155_c58b_6fd8;

        #200;
        key = 128'hbaa3_ea06_49b9_e42d_af80_6ff4_0b55_1de4;
        state = 128'hc4ec_2864_20d4_266f_80cc_b722_8a88_d693;

        #200;
        key = 128'h6287_54e0_91d8_8d27_26b3_6e45_2634_5a4a;
        state = 128'h9105_631a_78b7_1806_b5f3_c069_17d8_a347;

        #200;
        key = 128'h6000_0a59_5c86_2614_8a3b_d822_0daf_ce50;
        state = 128'h228f_2d37_63be_2cb6_3397_a735_8d6d_3ae8;

        #200;
        key = 128'he96a_b812_aa1e_3858_7426_b0e8_d51f_15fc;
        state = 128'h5a4d_cb53_c1a8_1e9f_5d19_f407_f13b_1966;

        #200;
        key = 128'h95d2_0f9a_21f1_fce3_d887_077c_aea5_1acf;
        state = 128'hfb68_76c9_6e71_8ff1_7394_467e_2f44_e560;

        #200;
        key = 128'h20a0_c011_d147_4fc7_d7d1_c3df_3ab8_9ed4;
        state = 128'h5877_2ebb_18c3_9a71_3aa8_213f_0474_e583;

        #200;
        key = 128'hd6b7_433c_5a79_109d_2e45_f179_b0a5_2ea2;
        state = 128'h2995_c7da_7470_d8dc_b601_627c_7a84_5d3a;

        #200;
        key = 128'h8ceb_85b4_8fdd_5db9_153f_6651_6073_1a72;
        state = 128'h3e80_b03c_35b4_079c_16ff_8c9f_d1a7_7084;

        #200;
        key = 128'h45cc_3c00_ac75_5368_047c_9bfe_7eeb_856d;
        state = 128'h6f20_18e3_0528_50ca_eaf0_47c2_1005_733c;

        #200;
        key = 128'h8c58_dbe7_72f5_10a5_c91f_eae4_e2a4_820b;
        state = 128'h55bf_a1d4_ab32_5b19_14cd_cda8_361b_db18;

        #200;
        key = 128'h4109_7e7b_b9f2_6fb4_210a_d53d_9596_a7c2;
        state = 128'hd0de_8df7_1e5a_c5f9_20ea_07e4_f919_aad1;

        #200;
        key = 128'h6463_a395_7bb7_907c_6537_8b00_fc27_076f;
        state = 128'hcefd_c6a0_3748_a653_dd61_2378_b719_580d;

        #200;
        key = 128'hf886_d5d9_2d33_b481_bfd6_e532_6f82_db8d;
        state = 128'ha322_332d_cca3_12fc_3f32_2627_ace8_3a71;

        #200;
        key = 128'hebab_91f8_afdf_0c4d_5ec0_be04_7299_dfde;
        state = 128'h4b65_e105_54cc_bf76_9046_d90f_aa83_b39c;

        #200;
        key = 128'h7b68_81eb_d661_2c88_6715_bb62_337c_ba67;
        state = 128'h69a3_1539_b4ae_3978_d55b_0c83_17eb_32e6;

        #200;
        key = 128'hf072_5311_837c_e4db_956e_8ca3_c3d2_2387;
        state = 128'h6f45_280d_86d5_f9c7_4e1e_e6cb_3795_1371;

        #200;
        key = 128'hf03a_b01e_d840_b3cb_55b1_2b00_a682_8087;
        state = 128'h255c_dd0b_2bf5_faaf_177a_163e_9054_f4d0;

        #200;
        key = 128'h50ba_bbbe_4286_9002_7857_e1ae_dc35_b4f5;
        state = 128'h3cb3_54ca_6c40_c097_ccb6_8976_f565_a714;

        #200;
        key = 128'h187f_c4db_fb63_2f16_bc05_bfa3_8494_2939;
        state = 128'h44a7_8947_b5c0_c97a_3aa0_9a8d_8b5f_668e;

        #200;
        key = 128'h6118_bd58_0437_24bf_3486_3753_918c_abad;
        state = 128'hdb8f_48c5_3e1d_fc63_0a8b_bbcb_7415_232c;

        #200;
        key = 128'h18b0_6e9c_322c_dd4d_3d55_b8f4_72e3_d40f;
        state = 128'h9bdd_39b2_8ce4_add1_ff83_7a27_7dc7_11b0;

        #200;
        key = 128'hdc51_574a_0d05_30c3_f4e8_ea1d_8f2f_0cfa;
        state = 128'h3d4e_6db2_91a5_9c8d_08c3_8b9a_1032_75a7;

        #200;
        key = 128'h7d56_f0cc_135d_0fe5_5180_1da1_3b9d_7d43;
        state = 128'hdddf_4243_8ccc_cd47_9e48_77ac_1e30_81eb;

        #200;
        key = 128'h356d_97a4_1298_cbfc_93e0_311d_419d_710c;
        state = 128'h1d0f_69a3_64a9_138a_4e32_4284_b9a7_f6af;

        #200;
        key = 128'hdb7a_9365_f468_34ed_c81f_535a_a944_8402;
        state = 128'hba95_749c_b409_c7c2_b482_bec0_3d20_5763;

        #200;
        key = 128'h2d31_a386_0942_2e4c_57df_54d7_c262_accc;
        state = 128'h95c7_3ba5_ab0a_4f4c_5d38_15ff_85aa_be63;

        #200;
        key = 128'h4432_6523_200f_338b_a2b5_ff84_35e4_b724;
        state = 128'h91a1_e40a_6e20_540a_b01c_4316_9031_0487;

        #200;
        key = 128'h92ea_8d4a_5463_9823_d89c_b8a7_ed12_3a93;
        state = 128'hf643_26a0_b0ec_48c4_e27d_1f2a_7844_3e17;

        #200;
        key = 128'hf399_9d7a_6c98_7c0f_93c6_0d96_b790_b487;
        state = 128'h8ce1_2ae1_35f0_09e2_b7ed_559a_5609_a1a8;

        #200;
        key = 128'he318_b9e1_4a9c_ec77_8e07_1eb1_2942_58c5;
        state = 128'hacdf_f0a7_6237_6dbe_f05c_4d0c_336a_9a43;

        #200;
        key = 128'ha7dc_9e8b_5013_15fc_fdb1_dbc3_c6dd_ab3f;
        state = 128'h4994_c4ac_87e4_d33c_807a_c4dd_1fad_0e8c;

        #200;
        key = 128'haa6b_9c14_2244_d9da_476f_aa54_7e6e_bf27;
        state = 128'h77bc_aa11_bfca_2026_a89b_a04b_44e6_3ff9;

        #200;
        key = 128'h8aa8_7ee0_6dd8_af93_d741_29be_083e_11fc;
        state = 128'h5806_5330_f6d4_d3d7_26ba_5127_55bc_feab;

        #200;
        key = 128'h4df3_2a64_cd4b_fcf3_f216_27f4_e012_2e8e;
        state = 128'h27b6_2a34_78d4_18e5_524b_4e31_47dc_f5c6;

        #200;
        key = 128'hf7ea_2f50_8bc2_fdb7_0f2a_4b1e_f6ba_cd9b;
        state = 128'hb84e_871d_d150_f579_1486_bd87_f929_c35a;

        #200;
        key = 128'hdff8_e612_07c8_da65_f778_f168_b06b_fbb9;
        state = 128'hdf23_02dc_0d55_921c_d44d_8c6b_b8f3_6b97;

        #200;
        key = 128'h9cfc_f467_973a_a773_f2ea_38cf_f51b_6628;
        state = 128'h49a5_60ae_f02a_07eb_9208_eb30_f3cc_9ba8;

        #200;
        key = 128'hfd75_a595_feeb_bea7_16a7_9d7f_e1a6_6a13;
        state = 128'hcd06_1770_f46d_1832_92d3_f438_e3e4_8ebb;

        #200;
        key = 128'h14f0_371b_9785_63b5_9bb0_5486_39b8_44c2;
        state = 128'h6622_08f5_6a46_ea87_4a41_f2f2_de2b_15f8;

        #200;
        key = 128'h7da6_5a5a_fa17_8b57_b4df_ee8e_7ae6_1b4f;
        state = 128'hc2ee_6fb8_6142_dd1b_e2b7_40ff_9ec0_2266;

        #200;
        key = 128'h4d79_ef21_816d_f9b3_4481_b320_bcf6_3c26;
        state = 128'h7133_668b_8e70_da56_983d_6a29_cfe3_c27c;

        #200;
        key = 128'h7c25_78a5_a9be_3c50_7f6b_7dbc_4a62_a237;
        state = 128'h58b1_f06c_0531_6cd6_6488_5008_04ca_fc29;

        #200;
        key = 128'h8aac_9c64_a5c2_1ad9_fade_b4ce_eddc_ae63;
        state = 128'h268c_11c8_ea1c_48b6_846d_5269_c9e5_ccba;

        #200;
        key = 128'h7d50_7aa6_fad3_8dad_451e_3a50_54c2_4bfa;
        state = 128'h3327_3fa3_fb94_6865_fa7b_c1f2_d703_e2bb;

        #200;
        key = 128'hade8_2574_ee1b_5827_8ca3_dc19_5688_d6dc;
        state = 128'h78b8_0633_9262_0823_0cf2_ed3a_0d7c_5482;

        #200;
        key = 128'h90aa_c191_ea75_1d30_affb_e3d7_6e4a_d514;
        state = 128'hd3f1_f2e3_6f27_fbd4_137c_1135_4c94_d36e;

        #200;
        key = 128'h26e4_57c6_6f1a_face_c229_4118_13f1_d1c6;
        state = 128'hba4b_af82_aa0b_f0fd_d31f_7fc4_0c82_155a;

        #200;
        key = 128'h40ee_234b_9302_77c1_48a7_06b4_e6da_65f7;
        state = 128'hda98_a66e_1366_b727_2bbf_69f9_8e2d_2ec6;

        #200;
        key = 128'hcda1_0f4e_78e7_e714_3521_951c_dd72_7cdc;
        state = 128'hcbf3_eac5_6ecb_99b4_0dbf_225d_0b1e_09a0;

        #200;
        key = 128'h747c_84e3_ec5e_3ef6_080b_64b0_98c5_3a49;
        state = 128'ha3b0_7103_87df_f29e_6ca6_cf86_cc62_4018;

        #200;
        key = 128'h2bc4_9ac1_c1ae_97b2_9419_6862_2b5a_54ac;
        state = 128'h75e6_8539_fdf8_3a14_6d95_c747_fa6c_26f9;

        #200;
        key = 128'h4664_f851_ea16_6044_7d5a_2310_d802_b45d;
        state = 128'hdd99_2c5a_76b3_9d73_6911_effb_27c2_5046;

        #200;
        key = 128'h0207_418b_fabe_6b3b_3d67_512a_ed47_3450;
        state = 128'hb6d8_3a3c_66bb_0366_28be_85ac_0a6f_89a3;

        #200;
        key = 128'h17e5_62f9_d189_72ce_3058_1063_cc0d_eecd;
        state = 128'hd829_56bf_c7f3_4f43_2559_ae91_7e46_9a7a;

        #200;
        key = 128'h16ee_0f40_6072_56de_667a_8e51_b679_ae74;
        state = 128'h6aa9_3b2d_93cf_4e40_cac5_fc64_fcda_dc05;

        #200;
        key = 128'h9514_e512_2583_3ad2_92d2_de19_a8ae_281c;
        state = 128'hee2e_bc40_60af_eae2_e46e_4a7b_ca27_b4f7;

        #200;
        key = 128'he2b3_a4ec_9621_3b33_98e2_e1a9_57af_140d;
        state = 128'h5774_e784_af06_20da_90a2_6147_2d55_3b7f;

        #200;
        key = 128'hb823_9008_7201_f87e_6da0_f274_ddb5_bd83;
        state = 128'hb9bc_f99f_1f71_802c_1c59_ad16_c410_195c;

        #200;
        key = 128'h00dd_995b_6eed_9446_a8e0_5c2a_852b_722b;
        state = 128'h20b6_8591_db9a_4731_40ec_2088_13b9_6da7;

        #200;
        key = 128'hf383_510a_30a2_b78a_bd61_8c61_0841_4df2;
        state = 128'h48f2_cc2e_d0a6_8a20_98fd_8d86_0a47_b487;

        #200;
        key = 128'hd801_8bc2_bce1_cef4_a5f5_50e1_80c0_0b3d;
        state = 128'hacb3_d72f_497e_846a_c85c_e0d9_9466_ed41;

        #200;
        key = 128'h3946_b43c_3a3d_066b_4f32_f624_5f33_a3be;
        state = 128'h5032_4b81_a80a_0e9b_1113_3c32_0397_e245;

        #200;
        key = 128'h515f_bef7_c235_c10d_0eed_8c8c_26d0_0c30;
        state = 128'h6e10_a336_2da5_b6c1_6469_a924_c6d9_f49b;

        #200;
        key = 128'h68aa_db55_2993_0172_950a_6acc_555d_7e8e;
        state = 128'ha6b7_6295_0c6c_5534_eb4a_d9f8_dbb0_8003;

        #200;
        key = 128'h9230_c54b_ba56_76b5_5582_5db7_2ee7_c8a1;
        state = 128'h0ca8_910a_f672_f0db_88e1_f8a3_5ef9_ead2;

        #200;
        key = 128'h46af_2795_7feb_d9c8_c125_7357_3d51_7e87;
        state = 128'hcca4_42a0_02d6_d98b_1d92_2be0_6143_d52a;

        #200;
        key = 128'h3bd9_a905_b605_f3ec_c758_213f_e611_9464;
        state = 128'hd00d_f89c_8008_0372_868b_7d41_9a62_84e8;

        #200;
        key = 128'h03f7_ae96_6af0_dcc4_e54c_6bc1_28d7_9424;
        state = 128'ha880_b117_376c_ef37_9755_4612_bddb_c66e;

        #200;
        key = 128'hf9c6_19f6_7a58_98ff_fb82_db84_2719_116f;
        state = 128'hc863_7a3e_12cd_cfb4_6194_7a90_d7ce_3c07;

        #200;
        key = 128'h1129_4dee_7cec_41d6_f062_c477_65f0_91f2;
        state = 128'h7cdf_cb64_8fe3_bb39_70f5_bdab_c21e_01c7;

        #200;
        key = 128'had5d_7ed1_c202_7f88_2f82_08e3_c679_c064;
        state = 128'h475f_9c15_e2ad_e91b_92b0_0eff_33e4_a455;

        #200;
        key = 128'h36c1_fb63_a64f_0eb9_694c_0e3e_ba98_4939;
        state = 128'hae31_6579_c0bd_ccc6_e01b_69c4_2e78_9ab8;

        #200;
        key = 128'hf231_5804_f01a_98c4_e6f7_77ac_8a44_8f83;
        state = 128'h2752_811f_ffa5_1bdb_5980_ff16_a694_5326;

        #200;
        key = 128'h391d_7ab7_d931_8ca0_8614_c042_69c2_3cd9;
        state = 128'hc8c1_26fa_43e3_bb70_3a60_c03b_e241_4dab;

        #200;
        key = 128'h08c4_2561_e27a_0ad8_d4f6_ac7d_866f_c72a;
        state = 128'h8d99_7c4d_e311_c327_a8de_ab6e_696c_1e9a;

        #200;
        key = 128'h8fa1_ecd1_83df_9733_b74c_a13e_2a0b_a7fb;
        state = 128'hb57a_0e39_442f_d56d_4018_e7e4_f94c_4867;

        #200;
        key = 128'hb768_f6f2_ef8f_40e7_ce68_e520_11fb_27cd;
        state = 128'h212b_2b99_8e78_bbf1_67ad_e7ef_dbfa_3da8;

        #200;
        key = 128'h9004_a419_7ad9_2b05_4d4d_65dd_0122_a96b;
        state = 128'h36d8_d8aa_103c_e5bc_4f89_8e40_1056_c08b;

        #200;
        key = 128'h6c42_f22c_c866_a1c9_6c79_32bc_f9af_d1c2;
        state = 128'h3013_36dd_cfa8_cb9f_b03f_4530_cec1_c7ef;

        #200;
        key = 128'hc1cc_f1d4_e967_eb58_04e5_0353_c77b_b755;
        state = 128'hd752_8647_c5fd_2a26_6a77_b653_5b3c_8d31;

        #200;
        key = 128'h4443_4345_bf2b_0c0c_f498_91e7_0860_ed12;
        state = 128'h630a_15db_c6ef_b17f_51fb_586c_c461_c209;

        #200;
        key = 128'h80b1_5ce1_966b_ac62_8f59_99de_d448_d6f4;
        state = 128'h402f_75f1_e79f_5a79_b83d_f1b6_e369_93cd;

        #200;
        key = 128'h28c1_6295_86f7_ca9c_5991_4512_642d_de74;
        state = 128'h1617_26d1_47c6_4b66_530a_3c7d_f296_a558;

        #200;
        key = 128'h60bf_9551_ebc0_20c6_7c0f_34c7_5d39_e70f;
        state = 128'h9c91_2d4f_50be_650a_1f8c_88da_4f4b_018b;

        #200;
        key = 128'h9c96_c313_e028_0d47_4d66_ad4f_1a38_e56e;
        state = 128'ha59c_6da4_b807_99ec_8d39_f0cd_f53a_75e7;

        #200;
        key = 128'h0689_f6b6_07b2_15dd_ecfd_99eb_9b7d_fad9;
        state = 128'h8d6d_cf0c_00d0_5619_1f32_b90b_0aeb_a655;

        #200;
        key = 128'h6066_7d7f_43fc_aace_30af_b0b1_e28c_f32b;
        state = 128'h8656_702a_3e6f_b2a3_2009_1db5_1ce0_0653;

        #200;
        key = 128'h973d_48ef_777b_0c7a_b871_3d06_475d_42d8;
        state = 128'h2f8a_981b_b12b_803d_0212_49b8_d026_93e9;

        #200;
        key = 128'h932c_6c72_4994_262a_17cb_f203_7391_37e4;
        state = 128'hf074_8662_e305_a566_d2c4_670f_8aca_869d;

        #200;
        key = 128'h377b_93a8_c43f_12bb_c5b3_459d_fc5d_1232;
        state = 128'h5926_c4ca_0e32_7f6b_e370_b242_693f_10b1;

        #200;
        key = 128'hc6f9_71eb_3e8d_5d33_6975_d1d3_4d1f_b5b1;
        state = 128'h72e6_1906_6ef4_5e64_82df_6eba_da0b_2cb5;

        #200;
        key = 128'h99e2_c964_b47f_76fd_7ab8_7da9_490c_aa5c;
        state = 128'h79a0_a6df_0668_ce36_ebf2_26d7_d093_a8bc;

        #200;
        key = 128'h25c0_6b94_08f1_5419_7d52_4d33_a45b_53d5;
        state = 128'h1533_1bd3_a4bb_01ce_87ae_7acf_375c_3deb;

        #200;
        key = 128'h4ff9_3982_0614_0a15_f531_100a_d6e7_9943;
        state = 128'h3575_d15a_7ea2_2b2f_1178_d3e5_044a_d057;

        #200;
        key = 128'h8891_e105_f204_a7d8_c2f0_c123_3e85_b5c6;
        state = 128'hc317_b2b2_ff7b_41cc_c734_b66c_aacb_9704;

        #200;
        key = 128'h69b5_c2db_690c_5914_bad1_daab_83ab_521e;
        state = 128'h8524_0c1a_1c96_6eba_9b35_7dba_d53c_1c22;

        #200;
        key = 128'h7630_dc55_6aec_939b_ec5f_92e3_8256_b2fb;
        state = 128'h0537_9703_24eb_cc8f_2712_58a2_412c_3e23;

        #200;
        key = 128'hbb0f_76d0_054b_9180_1cf9_f909_6326_6bbc;
        state = 128'h6adf_215e_4ede_98e1_b950_82a9_cd05_0224;

        #200;
        key = 128'h758a_821a_65ed_6caf_9758_65e2_576e_ad02;
        state = 128'hade1_7c0a_dd3d_25a2_c212_ad42_f092_d625;

        #200;
        key = 128'h35f0_8670_f155_97d8_6c01_9b46_2a4c_ce3c;
        state = 128'hc0d2_e51a_2f89_6c57_fc04_2d75_9566_453c;

        #200;
        key = 128'h05e6_7339_c336_f1b0_8d0a_22a9_0d8b_46fc;
        state = 128'h88e3_6ec3_d44d_c259_6214_d05a_c2c7_2ba8;

        #200;
        key = 128'h4a80_305a_430e_9b98_c211_3f85_5ddd_7f44;
        state = 128'h899d_33d8_b325_627a_5bac_bae4_73cd_9960;

        #200;
        key = 128'hcf95_3d82_f9b1_f455_6695_a6a5_06fb_59d7;
        state = 128'h7fb4_72cd_a5f7_acb4_2d3e_eaf6_bd32_159e;

        #200;
        key = 128'hd110_ddc9_113f_22db_d426_6657_9bda_b033;
        state = 128'hfc59_e025_72e9_8c07_11ff_1568_6a1f_cf75;

        #200;
        key = 128'hab7c_8eb4_fc78_7353_a080_710f_5b0d_8f8d;
        state = 128'h0c55_78b9_214b_69b2_1149_f5fd_9738_84f0;

        #200;
        key = 128'hb4bd_b0b4_53ee_c6fd_7708_6635_fc0c_2433;
        state = 128'h5af1_25c8_eaa3_bdae_7a0c_876c_dfd3_c534;

        #200;
        key = 128'h36ca_cf1e_9829_d627_7fac_8305_b193_27de;
        state = 128'h31a3_66ae_6d46_e935_f089_dc8c_7a5c_355f;

        #200;
        key = 128'h121b_ed8f_469a_ab24_66e1_9ae8_e716_1dcd;
        state = 128'h829f_3ad1_32fe_5f1a_a2a0_657b_0de1_e3cc;

        #200;
        key = 128'hace2_b33e_89bb_d2a7_0e48_0b66_72c0_e7fc;
        state = 128'hba32_5dbe_21d3_0bed_120e_e380_974f_d0b9;

        #200;
        key = 128'hd537_3cd8_8e38_aea8_1dd7_dd4c_72be_6817;
        state = 128'h0508_e877_d41c_e405_1510_be3b_18d2_43f4;

        #200;
        key = 128'hf36a_92b9_d464_c5f5_bac2_410a_ea15_14ee;
        state = 128'h8ae8_a657_7d62_1e62_7734_ae72_ef3d_d96c;

        #200;
        key = 128'hdbda_9e2f_64ee_c0ba_81b2_792f_c0fb_b878;
        state = 128'hbdc0_166b_b3b5_a902_2e85_563e_a83b_3a1d;

        #200;
        key = 128'h5b80_bd5d_ea96_747a_fcdb_2d26_51c3_00bc;
        state = 128'h4feb_eede_31ec_73f6_2f21_5966_9aab_ff94;

        #200;
        key = 128'h0a39_9c49_3c3a_a881_e646_69c3_6ec8_dd9b;
        state = 128'ha662_4f89_0aeb_5398_eb6e_e9e6_1f16_597f;

        #200;
        key = 128'h05dc_7f67_60c5_7cba_7c1c_2cf5_b2b5_ef6e;
        state = 128'h572b_ba30_fc8e_96c5_d7b5_1ccb_9480_5b41;

        #200;
        key = 128'h510a_31f2_1ed6_e0a6_a9c2_2547_ca8b_45a7;
        state = 128'h0e1f_add9_1373_1c8f_e39b_6ce5_863f_4e96;

        #200;
        key = 128'h7795_41e0_b22b_7ed4_7b90_263e_9ac4_f9e5;
        state = 128'h1b0d_66ad_2627_f921_9789_b792_4010_412e;

        #200;
        key = 128'h366b_a1aa_1178_7568_52a1_15d3_5cb5_8eda;
        state = 128'h09e7_be15_e948_2734_d191_d62e_7345_a841;

        #200;
        key = 128'h24c3_72b1_f6eb_e053_44a3_5b8c_34ae_d019;
        state = 128'hb13e_56ea_055a_7b2c_e722_c658_f7d5_361f;

        #200;
        key = 128'hf442_4eac_9725_5e49_f6c8_66a3_fa4e_0880;
        state = 128'h89e7_caa5_dd93_21ae_2feb_74c5_6942_89e7;

        #200;
        key = 128'h7c40_3490_50c0_83bc_16ea_31da_4ae2_fb7a;
        state = 128'h7c22_7e64_3bd8_15df_d0e8_cc90_d499_5b38;

        #200;
        key = 128'he8b4_47a4_e8a9_2e63_2944_0c76_ffb1_8a9b;
        state = 128'h0948_3e8a_0298_5a53_eb1a_4b13_cd04_2e94;

        #200;
        key = 128'h9baa_460a_4a6c_092e_8586_3a72_0e1e_6b8e;
        state = 128'h823a_2226_0845_e1cf_2729_dcc0_6972_91ad;

        #200;
        key = 128'h6bdc_a879_03de_8d3c_3c36_38e1_563b_3756;
        state = 128'haeae_1972_fe6b_387d_188c_5297_95b7_3ce4;

        #200;
        key = 128'h9f13_06ee_2d96_7f14_74aa_d1db_3372_9df8;
        state = 128'h867a_9e52_21e4_6fb1_ee9e_0e6e_2791_b22c;

        #200;
        key = 128'hf219_a5b3_4102_b074_6022_fe20_b6ae_5430;
        state = 128'h6aa0_a760_4f40_b63d_1fd5_08c2_bdc1_e8ae;

        #200;
        key = 128'h61eb_6824_de60_3fdc_21ab_0f71_5e56_8ffb;
        state = 128'h61d2_c785_f494_dbc8_4a40_6986_b53c_a5b3;

        #200;
        key = 128'h6c1d_0829_8c0b_d4d8_4540_a70b_eaa4_0730;
        state = 128'hf439_b506_09e5_3a17_55d7_00e6_7846_9ebe;

        #200;
        key = 128'h2e84_38a7_2728_ae39_78de_dd36_a3f9_c747;
        state = 128'hd452_f7ee_ab12_4da7_319f_35b3_d72c_54be;

        #200;
        key = 128'h702a_2f38_a875_f2cf_2c8d_1910_b3b9_ce64;
        state = 128'h2789_72b2_2f68_0c10_ca15_8425_7437_b0f7;

        #200;
        key = 128'heca7_392e_a8d4_ba2a_f198_91a4_ab98_e86d;
        state = 128'h57b4_9a4b_93a4_612d_2e44_e6e7_e1d6_057a;

        #200;
        key = 128'h91b5_e011_7967_fb39_1852_878e_90db_a7c5;
        state = 128'h4a90_942d_57ca_1fc2_7435_6d2e_5e61_89c9;

        #200;
        key = 128'hd737_8abb_3277_9030_6d9e_f72b_fff0_d7af;
        state = 128'h1559_bf66_886d_6278_318b_17db_e762_97f3;

        #200;
        key = 128'h4abd_dee1_3efb_1633_b675_70b6_49ac_b5d9;
        state = 128'hd0a9_a57d_3675_646a_d9e8_fc55_1e3d_21b2;

        #200;
        key = 128'h74be_6504_a5b9_2c0d_cfa5_9807_e6f0_b60a;
        state = 128'h5726_4e31_24c5_ffec_e699_c132_79c1_13b1;

        #200;
        key = 128'hb088_dfd3_d414_91bb_1207_136c_cba4_f876;
        state = 128'h825e_24d7_60dc_178e_6578_5513_8d5e_6796;

        #200;
        key = 128'h35e0_28c9_1ab6_7e07_4ae0_f7dc_5d63_3215;
        state = 128'hb615_8b93_d312_89e2_43fd_c02d_47af_622f;

        #200;
        key = 128'h3aa7_f47f_b0bd_b4da_6fe0_ab76_5ceb_ffe6;
        state = 128'h649b_4fe5_3caf_c5ae_49aa_ceb9_e159_09ef;

        #200;
        key = 128'hd7b2_7342_ea83_cea1_476a_c41f_daa2_6585;
        state = 128'h7ddd_c4c5_0172_1466_2e21_b792_2a06_4089;

        #200;
        key = 128'haabf_b1a7_e8db_2086_1616_2c78_d4f5_29ff;
        state = 128'h05be_dea5_d3bb_0743_f286_852f_88be_c765;

        #200;
        key = 128'hd052_dc79_d424_ec56_dbac_eda8_1a66_e8a1;
        state = 128'hdc0a_874c_e0e4_f872_3d12_294b_08e0_bea7;

        #200;
        key = 128'h6cd9_543c_18bb_337d_8233_f094_7154_7728;
        state = 128'h88d4_47bf_c6e0_c6c4_56eb_8e62_a03e_2049;

        #200;
        key = 128'h3c5a_dbe1_710a_57d1_7c10_0481_5458_3e10;
        state = 128'h692c_a528_6542_17d0_2231_0631_c647_fa8b;

        #200;
        key = 128'hcc63_2693_815a_ada7_9dc4_dd75_1aca_e73e;
        state = 128'hcc09_4b48_f0f2_d261_407d_3d15_f702_6532;

        #200;
        key = 128'h6135_80c7_bcd1_3fb6_1b2c_d548_047e_ec56;
        state = 128'hd99d_a66d_2e0f_198f_5259_428f_7f80_e1d6;

        #200;
        key = 128'h4c1d_0c50_ba93_040f_9878_2862_645e_fe1a;
        state = 128'h10c7_a626_4a4a_a71c_7beb_c869_b6c0_2b59;

        #200;
        key = 128'h38ea_8544_a1cb_23c0_d80f_14ff_f83b_d646;
        state = 128'h0b5f_f73b_faf6_cb99_f38c_a6c6_0687_f10a;

        #200;
        key = 128'h0c16_4cd7_95c7_3a5b_07d0_348a_c13a_9d12;
        state = 128'h18cb_be52_fd0d_b787_3244_bffb_366a_9fa8;

        #200;
        key = 128'haf83_9eb5_392f_a21a_49e0_1308_d558_3bb2;
        state = 128'h35ea_bd10_d20a_263e_ed4c_4fc9_13ff_1dc6;

        #200;
        key = 128'h1818_f42b_60a2_2cec_b08e_b904_13f8_03f3;
        state = 128'hf953_9d88_4ae2_14ae_e371_9120_778f_ba88;

        #200;
        key = 128'h7f78_d4a8_f804_47c8_1bc5_fa3b_bee3_c465;
        state = 128'hcfd5_ef7a_4152_c711_d972_745b_4663_ef83;

        #200;
        key = 128'h8fdf_810e_4d00_7ef1_3358_1f96_ca94_c1fd;
        state = 128'h1c1b_debe_93be_97f0_a26b_63c6_4380_f42f;

        #200;
        key = 128'hfc00_fa73_7972_5fab_27bc_6093_4599_f05d;
        state = 128'h4525_3023_54c7_5995_85b8_6ce0_5e70_0ce8;

        #200;
        key = 128'h864c_6710_235a_7416_6cee_e3f9_88cf_c1fc;
        state = 128'hc371_41df_d46b_5253_d095_02a5_f5fb_e321;

        #200;
        key = 128'h007a_fb41_6831_e5a4_90f7_84d5_9bf6_323f;
        state = 128'hcb69_50f8_a2c0_c5d4_2ff0_c738_89e1_e69b;

        #200;
        key = 128'haed3_9964_6cb6_30b7_7b70_02b1_e8f6_b095;
        state = 128'h641e_83ce_1111_41ec_6be7_bc82_278a_6df0;

        #200;
        key = 128'h0295_e624_36eb_0ed6_70cf_a87a_4087_d15f;
        state = 128'h31b6_d7e7_ddc6_f75a_72e4_dc86_f774_390d;

        #200;
        key = 128'h135b_01ee_91c0_15b4_82c5_36b7_db51_eac6;
        state = 128'ha2ca_b667_5df3_818a_b227_2bd1_2895_9161;

        #200;
        key = 128'hc0de_b0f7_0918_866c_b8ca_1991_f545_cfa2;
        state = 128'h1e1a_cddd_793b_d6b7_03c8_7893_46db_567f;

        #200;
        key = 128'h1bca_e208_1b3d_6fb4_02b1_1f55_6b92_7bb3;
        state = 128'hb644_347a_bdc4_3feb_ebda_dd6c_cc5c_638f;

        #200;
        key = 128'h3f7a_b045_5a74_8309_c618_bfd0_02e8_0684;
        state = 128'h15e2_6900_bc2f_d960_247b_11b1_fb1a_343d;

        #200;
        key = 128'hd875_343d_68e3_3955_4c17_7721_73fd_46f6;
        state = 128'h9053_d1ee_3aa1_e8db_e48c_1a73_ce57_820e;

        #200;
        key = 128'hda1b_9566_0ff3_6ec4_630f_4a19_c3e7_d028;
        state = 128'hcc9f_0017_c9c5_1739_aa3c_941d_ba2e_4564;

        #200;
        key = 128'h5d34_624b_1704_edb3_550b_4f3d_44a2_745e;
        state = 128'h8d70_22b1_cce9_2072_8fa0_dd93_a569_8b71;

        #200;
        key = 128'h9c39_6921_1f10_70cd_1d57_5882_f43f_5a48;
        state = 128'h08c2_7004_6a16_cc71_df2c_77ad_b9ec_7f24;

        #200;
        key = 128'h1d27_a72a_186d_c7b4_6d7e_0a6f_3a19_8371;
        state = 128'h9463_ffc1_fcef_aea8_0401_50fc_e2e4_9185;

        #200;
        key = 128'hb297_1c02_5289_55bb_a0bf_72be_a8d6_0146;
        state = 128'hdbcb_e127_c41c_cd83_9c32_8cd1_1457_cd55;

        #200;
        key = 128'h054d_7126_2994_1250_e3b6_1d67_ac79_45db;
        state = 128'hd67f_bd37_55b0_e16b_3ee0_fb58_3d2e_1afc;

        #200;
        key = 128'h3ff7_4a99_5388_e9da_5b54_b829_c6a0_f574;
        state = 128'he2c1_ce72_8300_d48b_4c24_8d9c_012c_b60e;

        #200;
        key = 128'hd6e6_5f38_cd3c_43c2_6726_350e_75ce_8ffd;
        state = 128'hb5da_2661_8b32_bef7_3699_cbff_9523_6c2b;

        #200;
        key = 128'hb458_5d89_151e_de30_22e9_715b_7416_d0eb;
        state = 128'h17ac_f131_8e25_a640_b29d_9dd1_37e2_1f5e;

        #200;
        key = 128'hdef7_cbea_551a_659b_f9b6_34d6_a5dc_a5ba;
        state = 128'h6d5f_eca2_85a2_57d9_1106_0a07_e6d7_90d5;

        #200;
        key = 128'hd1c8_cd05_565a_0ea4_3019_319a_30f7_658d;
        state = 128'h7d69_9acb_6ae5_5e7a_6fad_1f22_38fa_5dc0;

        #200;
        key = 128'h18cb_04ff_9d77_dfb2_a251_6e4c_1d1d_7e9b;
        state = 128'h467d_e58e_8796_0e24_6116_b9d9_3fef_e79b;

        #200;
        key = 128'h5cde_83c3_30f7_4f41_21db_d13f_efb7_2561;
        state = 128'h7f9a_789f_1538_0606_be7b_efe8_a639_f2dd;

        #200;
        key = 128'h4d6f_d11b_2f57_ce45_7b1d_16ce_1a6c_b8c8;
        state = 128'h84c0_1164_79ea_a001_ef21_5a95_9582_0bd0;

        #200;
        key = 128'hacf2_2224_f820_97ef_560f_f607_e2fd_7160;
        state = 128'h31ac_932e_7afe_f1a9_3014_d23d_00d8_f2c0;

        #200;
        key = 128'hc651_3bf9_f0c5_55f2_da49_6f24_6dc9_d2e1;
        state = 128'h670f_e580_5724_55f6_ead3_1709_b38c_d578;

        #200;
        key = 128'h14fe_d170_2045_f71c_74fa_e522_cb86_55ad;
        state = 128'h0a17_b236_ff20_7145_4c64_c2ea_47e6_78f4;

        #200;
        key = 128'hbe53_fd10_9c09_f172_8e50_8c0d_c62b_eb50;
        state = 128'h2b1b_08a8_f062_5f7a_1322_b259_3d59_9321;

        #200;
        key = 128'h962e_2508_13ad_104f_1d74_830d_d78c_5259;
        state = 128'h3663_95dc_5736_17f3_3f48_75a4_ef5e_3022;

        #200;
        key = 128'h070f_99de_90c4_d2ba_0860_9eee_5acd_d277;
        state = 128'h38a1_44df_57d4_2e1b_cf9c_338e_0b41_0d1b;

        #200;
        key = 128'ha2fc_bdd3_57ed_5d1c_b9a6_6839_0eca_a73f;
        state = 128'h3632_3659_874f_752c_a0f7_cd1a_c2f4_852f;

        #200;
        key = 128'h2e18_8cca_1b37_757d_9773_e8b0_e4a0_07b7;
        state = 128'h63cf_97ec_28db_9c6f_973d_5ba0_d613_2793;

        #200;
        key = 128'h4558_496c_200e_83c0_c73f_5269_5cf9_3b4e;
        state = 128'hf6c0_afda_5b86_3a36_660d_50cd_e803_215e;

        #200;
        key = 128'h83d4_27be_bd21_5cc0_ae49_bc62_45eb_f084;
        state = 128'h5a98_5a37_dcc4_3ab0_c402_3e6c_e4c4_f292;

        #200;
        key = 128'h4c59_d358_fd98_6478_534b_79c1_8cc0_de23;
        state = 128'hbffb_c970_2d79_b6c2_7b36_675f_c66d_99b5;

        #200;
        key = 128'hdcc4_6d5c_4b2a_a19b_efd8_3544_c3cc_b857;
        state = 128'hcc13_960b_b860_ecef_883e_7566_c73b_3564;

        #200;
        key = 128'ha9a2_1287_219c_4ed2_56f6_32cc_a5b8_8a21;
        state = 128'h3a64_8016_d58f_df91_3a73_3ea9_acff_530e;

        #200;
        key = 128'h7aeb_1e81_1637_e01d_8378_9b87_0ec7_f6ba;
        state = 128'h4732_0f75_4af1_3ab6_4e1c_d8b7_3a59_3048;

        #200;
        key = 128'hcaa0_35ac_4eeb_bee2_4dc2_a8e7_9858_05c5;
        state = 128'h1ccf_0a3b_19a3_1a1d_54da_fddf_e30b_7a0c;

        #200;
        key = 128'hb2ba_337d_2ff2_4662_01ae_6d00_e810_c393;
        state = 128'h3b83_6d9e_a19f_e4a3_6deb_af39_be1c_f70a;

        #200;
        key = 128'h28c3_a70f_cbc4_000f_2840_2668_1b10_8bd0;
        state = 128'h44ca_d456_14b9_83d1_b2db_8db9_3bd6_3be4;

        #200;
        key = 128'h3ee3_9e73_74ee_4c59_e13e_09c3_a7ca_1cd3;
        state = 128'h220f_db80_f7b4_e244_c2d7_7785_a67c_24b3;

        #200;
        key = 128'h18ab_1ce7_5e16_309e_46be_8d53_400f_e6ab;
        state = 128'he1ca_4a06_9d02_9f7a_bc09_8d27_7bbc_ffb2;

        #200;
        key = 128'hc927_0d1d_4503_d883_81c9_2b70_dbc9_1122;
        state = 128'h2c07_6b80_94c1_1265_ff83_fe31_5539_dc86;

        #200;
        key = 128'h7069_4480_0682_2b3a_3a06_7e0d_7995_00f5;
        state = 128'hc039_9ae6_4849_a54e_d5ae_b574_3cd8_735f;

        #200;
        key = 128'h7fe2_4caf_6c44_d92b_a05d_913f_b53e_2991;
        state = 128'h3c5f_323f_fd20_71b1_32c6_b591_a164_87b6;

        #200;
        key = 128'h953a_4ef9_2b05_a18a_8c60_d7f9_f658_c3e4;
        state = 128'h5a5e_92ce_f234_5ad9_7dc1_ad9f_a91a_6e39;

        #200;
        key = 128'h0df3_60da_5392_3e94_1991_35d9_5210_84cb;
        state = 128'h6343_9311_e31d_9e07_79ff_2935_fbe6_617e;

        #200;
        key = 128'h19e8_81da_24e1_0158_f4ab_5c43_3836_6acf;
        state = 128'h315d_a7c8_172c_0718_028d_3a62_495e_b7f6;

        #200;
        key = 128'hcf52_4436_45c3_75ef_ccf5_27be_cf68_b693;
        state = 128'h8c37_b599_a4a2_51d5_715f_f821_d0da_3918;

        #200;
        key = 128'h300f_611f_7904_b5d2_fe48_d0ab_07d1_d24b;
        state = 128'hc5fd_146f_06aa_86e6_54b9_669b_fcc8_9d01;

        #200;
        key = 128'h047a_cf3d_f4c8_0b3c_6e1c_9d41_09fb_9c3e;
        state = 128'hb0c8_80cd_ed2a_dded_bf8d_0509_ecf0_4ff9;

        #200;
        key = 128'h0aad_6731_66f8_3d7f_9eb8_511f_e51f_6f6a;
        state = 128'ha014_f163_1da9_017f_53c6_383c_1d81_6d9f;

        #200;
        key = 128'hb3df_90bf_8373_a157_bdae_2285_a863_502d;
        state = 128'h8e44_a2b1_ee2f_5bd4_ec98_6c6d_c4d4_3146;

        #200;
        key = 128'h8b7c_a15a_e382_e6c8_5e37_4ffe_413e_6db7;
        state = 128'haa9c_240a_26b7_519a_2cd0_b235_606a_bf4b;

        #200;
        key = 128'hff48_c895_b408_8915_e10a_1de1_4c1c_a587;
        state = 128'hda45_b3b4_5853_c6b4_d1c2_b372_4e6c_8d16;

        #200;
        key = 128'h5c2a_dc62_6d87_9b23_2af0_1864_8520_fc33;
        state = 128'ha573_e770_10d6_2d7d_c400_0a1a_9163_9ee3;

        #200;
        key = 128'h9b48_6b29_030d_fa43_a6e0_bc64_ff90_3872;
        state = 128'hc0a4_b776_cf57_942e_c0ab_773e_cca6_1c9e;

        #200;
        key = 128'h6468_a5c7_3947_715c_a181_fe12_6127_7861;
        state = 128'he6c1_f772_d9be_4fb4_bc0f_65be_6579_1cf0;

        #200;
        key = 128'h08db_dc0a_8362_8082_aab8_bbda_d81b_af25;
        state = 128'h1f32_a4a4_1c88_e273_9d24_1248_2eec_f103;

        #200;
        key = 128'hf42d_bee5_c997_4e13_0f08_b7b8_7909_3494;
        state = 128'hf7ec_8ca7_b90a_d1e7_f46d_ef83_6deb_24d8;

        #200;
        key = 128'h8542_fe43_7f85_bfdc_e13b_fa6f_14bd_8d78;
        state = 128'h4507_e986_b8c5_67ab_f198_83db_bd12_dcda;

        #200;
        key = 128'h3ee7_bfdb_13bf_8015_9510_6695_5d1d_2be1;
        state = 128'h4f94_28b8_3c40_4a79_8c92_8e69_f485_4892;

        #200;
        key = 128'h44c9_0993_74dc_ba07_c692_6ff7_6c65_6efa;
        state = 128'h686a_17a2_3413_1331_d12d_f311_03fc_1637;

        #200;
        key = 128'h388c_0af4_d049_dedf_64c3_444a_ca4f_c703;
        state = 128'h4001_1851_6a49_23f8_546c_fbb1_e643_eedc;

        #200;
        key = 128'h819f_7f8d_456f_7b0b_8496_9d5b_60f1_9b76;
        state = 128'h1017_30b8_95c3_a822_05d9_cefa_5b42_9cfd;

        #200;
        key = 128'h2dad_74cd_6bb4_cb36_9b4d_220b_7170_a486;
        state = 128'h22b0_5047_8632_6c72_49ca_85d0_c6e3_aceb;

        #200;
        key = 128'h19fd_d3db_4e7c_1143_483b_0298_15f3_298d;
        state = 128'h489b_05a7_0bf3_6ed2_d028_b1b2_e5b4_6c9e;

        #200;
        key = 128'h1d40_c01d_ee25_086c_1cc6_0810_83e6_38fb;
        state = 128'hbb0b_345c_3b94_619c_57d7_b9e0_707e_739e;

        #200;
        key = 128'h645a_31e3_1ed7_bf4f_eb54_6291_928f_b264;
        state = 128'h7a3a_b12f_227e_1d44_a3a7_cad7_9308_425d;

        #200;
        key = 128'h77fa_4465_4cc3_1b8c_7607_c02b_132b_2d16;
        state = 128'h4adf_bbf4_c7ce_e093_32bc_243c_df82_37c5;

        #200;
        key = 128'hb7a6_281e_9e76_34ea_5176_5268_abb7_7f72;
        state = 128'hcd26_b855_878c_01bc_421a_f551_e075_5460;

        #200;
        key = 128'h83bb_b845_f526_7d34_dd35_27af_cd79_e0a4;
        state = 128'hfa92_cbe8_bfd4_0119_f476_80f6_b097_d28f;

        #200;
        key = 128'h6184_0741_572e_5d36_07c2_3757_7744_d085;
        state = 128'h89c1_0ef9_2666_51a3_c3f9_a041_10cc_14f7;

        #200;
        key = 128'h7568_b0f3_6f5d_e3fb_427f_8a33_aecc_5b1b;
        state = 128'h0551_c49b_3718_68ab_47dd_2300_68ca_ae73;

        #200;
        key = 128'hb1d3_cf0c_c516_668f_d589_c575_0025_6df9;
        state = 128'hf5b2_bcea_668d_0cc2_08f3_d2e7_169a_515a;

        #200;
        key = 128'h87d0_dcc2_7c0f_4415_9d5b_e9b1_7f2f_8583;
        state = 128'h43d2_c67e_bdaf_588e_ed49_e44f_0179_5a30;

        #200;
        key = 128'h8d2d_538b_280c_4816_d7d1_8fce_7002_be3a;
        state = 128'hb327_3b65_870e_802b_740d_1054_6f60_cfd5;

        #200;
        key = 128'h53f0_623a_7bbf_d3f5_e718_1acb_192b_f900;
        state = 128'h9936_cc69_a833_c4ac_cf4d_e8bc_3907_48f7;

        #200;
        key = 128'h9056_c5b1_0f70_b267_a297_2173_ca41_9de6;
        state = 128'h5d75_a134_1385_ff3f_7e94_ab35_1e85_53c4;

        #200;
        key = 128'h4c3e_cb55_05db_1dec_83d7_b09e_04dd_c99c;
        state = 128'he0b0_4518_3726_9664_d257_6c09_acc6_0cc4;

        #200;
        key = 128'h23ec_6dbf_7531_66ad_c899_533a_ff5e_217c;
        state = 128'h4e49_654d_326c_b821_dd6f_031a_966c_5358;

        #200;
        key = 128'hb446_63fb_2121_44d1_fcff_3317_acc6_f692;
        state = 128'hf741_0a2a_a4e2_524a_b574_9083_b87d_9a38;

        #200;
        key = 128'h859e_d828_724b_37cc_ee10_dd9d_3ec3_3992;
        state = 128'hfce3_a3e4_71f3_06a7_ba5a_f93d_1f14_c250;

        #200;
        key = 128'hbba9_ded3_515f_4353_64f2_dc84_f206_87e2;
        state = 128'h2cb0_8de5_2ef8_65a2_aab3_959b_89f8_ba44;

        #200;
        key = 128'he099_d449_ff46_0f54_3d51_7892_ced6_db4a;
        state = 128'h8ebd_3354_811e_316d_dcea_ea4a_9719_c56f;

        #200;
        key = 128'h1299_9884_f330_f725_e602_81c5_b777_da7d;
        state = 128'h9898_2964_1f25_ea05_8c80_068e_2379_e4df;

        #200;
        key = 128'h690e_cb17_a820_bc36_c60f_4606_8bb5_20dc;
        state = 128'he1df_5608_d8b6_5556_c928_6e71_1d90_88b1;

        #200;
        key = 128'h85af_ef5b_fd2d_8f1e_93be_8e6d_29b3_0e0a;
        state = 128'h00c6_6164_3dd8_0674_02e5_c3ec_6d89_4953;

        #200;
        key = 128'h65cd_8236_733c_cdb5_80af_95a4_4060_74c0;
        state = 128'hb667_9390_8dd8_75cc_720b_3f2a_172c_e3ae;

        #200;
        key = 128'hd912_ba7f_03ce_ce5b_80bf_ef03_1500_2f31;
        state = 128'had75_bd2f_2dc7_fad0_83a4_7f62_a96b_bd93;

        #200;
        key = 128'hca81_2b63_243c_612e_7c45_1817_224a_c4dd;
        state = 128'h5a7f_624c_e491_6978_3782_39db_a0d0_9f53;

        #200;
        key = 128'h7222_5541_2231_85a8_195c_d32f_8340_4937;
        state = 128'h6b16_4fcd_fa91_d171_b7af_f7ee_f53a_bf91;

        #200;
        key = 128'hd8c6_3a53_41a3_9a8d_9bd4_00f6_73c9_11ff;
        state = 128'h5d69_a564_b76e_9a32_42a1_9ee2_0321_31a1;

        #200;
        key = 128'h8b2f_0058_66fb_329e_5260_a501_45b5_b43a;
        state = 128'hb3af_06f0_5d97_bd85_395b_57a5_acb5_e4e4;

        #200;
        key = 128'h24d1_60b5_905b_b41a_92cb_36ad_ff4a_4e2d;
        state = 128'h614a_9d67_c390_5e8b_5004_45d1_faf5_05b1;

        #200;
        key = 128'hda38_8021_7a87_b126_9fde_796f_bb53_4b91;
        state = 128'h4bf3_ae62_63c1_2c06_42e6_2685_75b7_da73;

        #200;
        key = 128'h8667_1a48_a445_a5eb_45a5_8533_45a8_dd2f;
        state = 128'ha88c_0bda_d541_8b96_0ed3_11fe_931d_75fb;

        #200;
        key = 128'h0008_f422_2df0_ab27_5f5c_5237_d1da_92c8;
        state = 128'hc11f_b781_c47f_18b4_2a72_62e1_3c99_1208;

        #200;
        key = 128'h1c03_d2f7_d053_135b_2fca_0789_2b8f_c488;
        state = 128'hab2c_4454_5baa_a5b8_4beb_9274_6a0d_431a;

        #200;
        key = 128'hf47e_0327_d0df_8c71_4252_d986_8520_e0a7;
        state = 128'h08d8_5225_f8f1_7aad_c661_1ae2_0a6f_05e8;

        #200;
        key = 128'hc2df_744b_70dc_4d17_dcc6_9fc0_7be6_fc99;
        state = 128'hd8fe_18c0_684c_d353_d1e4_8674_7017_5439;

        #200;
        key = 128'hcee5_3c29_f5e5_241d_629a_6ee0_6266_3eba;
        state = 128'ha163_cf56_8e30_2f2f_b98d_f847_f2d2_0ef0;

        #200;
        key = 128'h22ba_2f99_55d7_6afe_9423_e037_4139_13ea;
        state = 128'h30da_5db0_427c_0f26_1955_1df0_8df1_dc70;

        #200;
        key = 128'h0a84_e72d_f1a0_0871_e9a5_de09_90ed_07c6;
        state = 128'hec61_af6e_4830_71c8_c087_5804_fc37_a4eb;

        #200;
        key = 128'hf751_11e1_f83d_9faf_a4d4_2276_0479_9a0b;
        state = 128'h0189_b682_3ee8_2bdf_0c9c_8427_a3ac_36d7;

        #200;
        key = 128'hd227_44d9_85af_51f9_bf29_555c_7e33_09d1;
        state = 128'hb74d_5e8f_a2a4_bc04_bcd4_ddaf_c7d9_522d;

        #200;
        key = 128'h7fff_89da_f1f7_3cad_2216_816e_59c6_f909;
        state = 128'hfadd_b7b7_d786_365f_bb2d_2421_7b8d_4f34;

        #200;
        key = 128'h45f5_aa7e_0d3c_2f6f_d488_8e60_6b1d_526c;
        state = 128'h8696_84f1_95f4_aa9c_40a8_beeb_60ee_c5dd;

        #200;
        key = 128'hfd19_8bf8_15ec_cfab_36cf_51e5_679c_b1ed;
        state = 128'h06f9_d945_bf5e_9d3c_f9ba_3ab9_3504_70a3;

        #200;
        key = 128'h255d_8a53_264d_e0cc_52ca_ae0d_5b9d_e3ab;
        state = 128'h698d_7a83_37f5_9d49_6d26_1d9d_bc95_1c80;

        #200;
        key = 128'hb138_d38f_5bd7_2eb3_1cea_9998_79fa_3840;
        state = 128'hc61b_03e0_d397_e6fc_bd76_d6cc_48fd_29b2;

        #200;
        key = 128'hc908_6275_e52c_c228_df8b_0232_8353_21f7;
        state = 128'hc006_7628_4ba8_e5c4_6407_2160_8300_5ce1;

        #200;
        key = 128'h1339_cc87_36ee_359c_2311_0388_e8e7_2b0c;
        state = 128'hd427_9dd6_3732_bbf8_dd16_73af_f82f_e205;

        #200;
        key = 128'h5524_5502_7235_7b89_4692_89e3_7a2f_8fad;
        state = 128'h0084_8e98_2778_cbc7_80ad_40c2_92e6_405e;

        #200;
        key = 128'hebef_854b_c520_8385_f73f_c11d_e314_645a;
        state = 128'h1908_8ce7_ddbf_48f9_1a4b_b918_de03_d320;

        #200;
        key = 128'h9c59_189a_791e_c325_ed9a_4ce5_1c0c_33db;
        state = 128'haef0_51b3_a1d7_db74_3840_ffa6_1ae3_6666;

        #200;
        key = 128'h750b_a003_4736_e6df_b327_164e_b6f9_11bf;
        state = 128'h40fa_fc9b_a4f8_6790_f9ad_83ac_45ec_fbe6;

        #200;
        key = 128'h5b44_f8e4_1d66_60d0_bad6_2081_23db_b3f7;
        state = 128'h757f_d30c_20da_1873_b108_7c3c_72ea_f123;

        #200;
        key = 128'hcf28_3ef8_59e0_abee_b925_6195_7e94_9648;
        state = 128'hb667_95b6_dbc6_44db_0416_45aa_0569_5b83;

        #200;
        key = 128'h0804_71ea_3037_533b_8ccd_90d1_c0f0_f9ed;
        state = 128'h6103_73c1_05aa_4dd5_acab_4d18_bb6b_6c45;

        #200;
        key = 128'h5355_9ae1_56f5_e98d_7bb2_afbe_af86_00f9;
        state = 128'hd33a_5567_818b_6f44_93ba_8a78_53a7_68f3;

        #200;
        key = 128'h2718_1ae8_5bc7_2ee4_87b3_7451_dc1c_7531;
        state = 128'h3d7b_e86e_db5b_032d_03fe_0b7f_955e_07cb;

        #200;
        key = 128'hb3d7_9317_c4ff_cd33_b16f_bb49_c761_98ed;
        state = 128'h05d6_f5eb_89c0_fff5_4bfc_88a8_c03b_9a05;

        #200;
        key = 128'hb440_ca31_4b52_9e31_2488_e41f_df83_8858;
        state = 128'h1eb1_00bf_8b84_7444_28fe_7e27_59f1_3748;

        #200;
        key = 128'h6941_a817_8dfa_d67a_c1e0_b46a_3806_8e1f;
        state = 128'h164c_d7d9_17af_514d_e158_2942_2b51_ca4d;

        #200;
        key = 128'hf6d4_c765_3a37_923c_8cec_f87b_972c_568c;
        state = 128'h06e5_f55a_8a5f_9f99_edac_6029_ef51_27a5;

        #200;
        key = 128'hbb48_4659_f756_443e_1e9c_9371_e45e_1ff3;
        state = 128'h25c4_72d5_1576_fd77_a8a9_07a7_08ba_68e4;

        #200;
        key = 128'h2ebb_ba44_532d_8fe1_e8c2_7324_0b8a_129e;
        state = 128'ha7b8_8205_8917_b291_ec3d_85ad_c9b3_5dd7;

        #200;
        key = 128'h2b6c_ebf0_e172_da7c_0fbe_0a2b_b8c7_f20e;
        state = 128'h61a1_8ccb_7f30_0c62_9473_f65b_72f2_1006;

        #200;
        key = 128'he900_1c88_8261_90c6_c37d_e438_7ac7_55b5;
        state = 128'h6c48_2931_9eeb_7207_f33e_293c_c0e2_4fca;

        #200;
        key = 128'h0935_6f3a_e384_3c7b_fc32_2f0d_2600_987a;
        state = 128'h9e61_ea00_f56f_46f3_90e9_5af0_1eea_510e;

        #200;
        key = 128'h4515_8f55_9938_dfea_b523_2014_5261_1588;
        state = 128'h5910_670a_3fc7_6823_c001_0f97_0f83_3ad6;

        #200;
        key = 128'h05a7_6a97_61ac_ff07_1aee_7ad1_eca2_97da;
        state = 128'h1d24_ce8d_f4f3_c429_e175_c612_37a6_dde1;

        #200;
        key = 128'hd662_3c67_d97b_a116_5dda_c685_f3a4_f7cc;
        state = 128'ha703_629f_993a_2466_8f0c_3190_a57e_ca1d;

        #200;
        key = 128'h6761_3da7_7edc_7d8b_1ffc_9ac0_0d66_57fb;
        state = 128'h02ca_bfaf_268e_0780_64fa_f9fc_1393_7532;

        #200;
        key = 128'h4ad0_0292_9415_b0de_bcfc_121c_57a3_6c44;
        state = 128'ha07f_d694_64e0_db80_ae0e_18a4_a141_ef17;

        #200;
        key = 128'h4eed_b235_695b_67c9_ca87_ee4f_ad99_f17a;
        state = 128'hca13_1bcd_df28_4857_a2d3_e0cb_3230_5b68;

        #200;
        key = 128'hf2c4_3a34_810c_ba05_7561_6bef_e8bd_fb0b;
        state = 128'hc919_5ae9_875f_a8ed_bc2c_96a3_6b45_4481;

        #200;
        key = 128'h0116_72aa_0110_3c83_acbb_2e8f_b40a_bf46;
        state = 128'h92eb_8002_ccae_b80b_07a5_07d4_a6a4_cace;

        #200;
        key = 128'hd618_645e_8879_bda0_2e8d_efde_7adf_0e09;
        state = 128'h37c5_7631_9390_2e13_3c3a_4ffb_ae24_ecd1;

        #200;
        key = 128'h8361_4756_5e35_a27d_e57c_87f0_8b99_c830;
        state = 128'h4ef6_6674_5844_f12f_01db_c532_a4cc_6e3a;

        #200;
        key = 128'hbde2_04f5_93af_3eba_eea3_3027_2f44_8622;
        state = 128'hc2d4_dd9f_933b_70f7_6eb4_9403_94df_0e90;

        #200;
        key = 128'h72ab_2b02_f077_0def_a40f_444c_dcb3_34b4;
        state = 128'h2967_b405_7538_6ae2_34c1_88c9_ef8f_c020;

        #200;
        key = 128'h95dd_0a0b_39e1_b348_c43d_fafc_78c0_0a10;
        state = 128'h3e90_6f86_3581_b634_5b07_c4aa_7879_34e5;

        #200;
        key = 128'hbb22_cb5e_53c1_b503_2bf9_efdd_3437_d17a;
        state = 128'h32d0_40be_6156_77d0_f92c_5cae_e935_27eb;

        #200;
        key = 128'h145c_7581_f6b8_1a41_0e3d_63a0_d414_5737;
        state = 128'h11cf_f29f_4f95_4ff1_66e5_eab0_fc7c_c661;

        #200;
        key = 128'h906b_13df_cc09_4c12_ea10_fb08_0d7b_2154;
        state = 128'h6fff_b739_9862_03cd_4ca1_6526_322c_cb83;

        #200;
        key = 128'ha2b1_4dce_f3a8_81f7_7cd5_654b_3e3f_5f3d;
        state = 128'h909b_b10c_c072_6af3_3d32_cd92_2238_7656;

        #200;
        key = 128'hc1a3_f3f8_1f82_78a2_69ed_fa1e_1dfe_e431;
        state = 128'h699e_32ba_185a_81a4_49b1_01eb_0cc5_1a8e;

        #200;
        key = 128'h7d55_47e5_336f_31d7_b34a_2199_3dce_fe1c;
        state = 128'h185a_d08d_17c9_9859_814d_7e59_15f2_56ac;

        #200;
        key = 128'h9a99_0c33_0d86_a097_72f5_32d3_6943_48c3;
        state = 128'h1b38_e7b6_5cfe_5b01_6f4f_fa6f_7275_7a18;

        #200;
        key = 128'hf9c4_ea08_c79a_4581_cc72_782d_2e02_54fe;
        state = 128'h2c3e_4fe1_dd99_4f47_3c75_97ae_28fa_967c;

        #200;
        key = 128'h4028_ef9a_0b35_acf8_dfa3_846c_031a_f47c;
        state = 128'h55aa_1d5c_4b73_a372_5c7e_f119_beb2_fd99;

        #200;
        key = 128'hd503_5714_0de2_13c1_2fb6_6281_7c07_8481;
        state = 128'h1aeb_2ac4_0303_7c09_33a4_882c_ad4c_b37f;

        #200;
        key = 128'he724_7f88_b167_92ff_ff29_c928_1ecb_0df1;
        state = 128'h3549_cfa7_89e7_a929_17bd_b3b0_5094_05cd;

        #200;
        key = 128'he02a_99a7_cb6e_2308_2ab4_b466_d18f_fbe6;
        state = 128'hce01_6b44_aee5_d35c_f1bd_5719_a01a_a02f;

        #200;
        key = 128'habbd_5acf_ae1a_8418_047e_c306_d68f_4611;
        state = 128'ha6cb_ec6c_53c9_0131_bbbb_7c8e_471d_92d8;

        #200;
        key = 128'hf2b7_73aa_9c92_a30b_288a_c85c_b780_5185;
        state = 128'hc6da_3905_d292_e493_fa8e_11e2_6ade_eb48;

        #200;
        key = 128'h48e0_b219_4d32_1db7_3acb_9db6_cfca_4a4a;
        state = 128'hb0de_60a7_2851_29c8_eb01_b60e_dcf5_c462;

        #200;
        key = 128'hf1bf_5732_3f72_0470_5419_4df2_4623_30b6;
        state = 128'hfdc9_bd19_6cb8_8ed7_ddd0_31e2_a571_6313;

        #200;
        key = 128'h4a0d_2a5a_26c1_3005_1a4f_c730_99b8_0e0d;
        state = 128'he92d_6cdb_6803_368f_c7f5_36d5_3dd8_1f46;

        #200;
        key = 128'h1ff0_6982_b4e7_3be3_5f13_7df0_11ff_150e;
        state = 128'hc0a4_f3ac_a6f0_4e09_e0b0_2b59_d134_35f0;

        #200;
        key = 128'h4f44_030a_7cec_08ec_a3e3_1957_a75e_6e6b;
        state = 128'hf1f3_ec0e_1d06_ddad_c5fb_28ba_bfb2_aff8;

        #200;
        key = 128'h679c_78d4_982f_f832_a3a7_dee4_56ff_ad14;
        state = 128'h14d6_03c2_8798_28ef_b9c5_d66b_b3df_2779;

        #200;
        key = 128'h91a0_1ebb_5e78_b949_cbea_5dba_aa97_b28a;
        state = 128'h1d8b_b133_64a4_08da_24d3_7d7b_22ce_509d;

        #200;
        key = 128'he7b1_6837_725f_95f6_0a80_8db1_0839_6f82;
        state = 128'h1414_7c45_4351_2584_cc01_7c41_5529_29a1;

        #200;
        key = 128'h4c13_df0a_c4c5_74e6_1682_1b82_ddac_020e;
        state = 128'h19e5_502f_660e_5fe2_13e6_1dd8_368b_160c;

        #200;
        key = 128'h7661_6694_712b_1f05_5179_c94a_9395_fba9;
        state = 128'h73f7_e358_26ec_b4b4_a369_7156_70cc_115a;

        #200;
        key = 128'h5963_4079_9ea7_f9ec_c1ec_d0b7_0088_73f3;
        state = 128'h510e_3fa0_edf0_f93b_da79_3f3b_c07b_50fa;

        #200;
        key = 128'hcc26_587d_cea2_7193_5823_216d_a241_dc43;
        state = 128'h541d_e7a7_8481_44d7_e855_cca0_ef9a_a5eb;

        #200;
        key = 128'h5596_fedc_7ab0_443e_1c1a_d821_0fce_2ac7;
        state = 128'h1039_6721_87b9_ba97_3bbf_6e57_8771_2ab0;

        #200;
        key = 128'h10eb_81ec_cc72_ffea_9375_1dff_a023_f329;
        state = 128'h61f5_8ebf_43cd_ed47_85fd_0d04_e3b6_d9d7;

        #200;
        key = 128'hb070_6985_0db3_9ac8_0a6b_daa6_bc6a_16f0;
        state = 128'h6298_75ce_a227_5eb9_49f1_522c_2a88_172e;

        #200;
        key = 128'h571b_a70e_42e7_ce67_f7cc_a0d1_3759_f636;
        state = 128'h7f6b_fcf4_2c77_4e96_8bfa_cd44_68f9_a0a6;

        #200;
        key = 128'h4c15_d21f_6639_72d2_1b04_9b78_8c47_808d;
        state = 128'hc6de_fda7_7ce8_fed6_fd6a_9c62_c80b_0339;

        #200;
        key = 128'h038b_01fe_f026_3eb2_b2c7_2339_c9dd_e67e;
        state = 128'hc788_26cb_b13e_af83_1520_ad83_1c97_3595;

        #200;
        key = 128'hea5a_dc46_a41d_5bf4_437c_125d_3572_2b1f;
        state = 128'hd9bc_0786_0ab3_005f_89c5_579f_6986_9931;

        #200;
        key = 128'heea5_1294_5f4a_bc95_e4fd_467c_7983_1232;
        state = 128'h1bd1_b4af_9ae5_1682_9ba0_ae19_1bc2_07ac;

        #200;
        key = 128'h3ed7_7605_1981_8c88_6100_6b4c_1bec_3ed1;
        state = 128'hcfc8_6c33_830c_bcb0_08f6_691b_ed4f_087b;

        #200;
        key = 128'h0848_e800_f670_3d86_050c_662f_53ea_a633;
        state = 128'hdf0e_7c3b_38ec_4c95_2a89_15ab_0843_9cde;

        #200;
        key = 128'heaa6_ec81_3896_1da4_e7d2_ebda_5f3f_86e0;
        state = 128'h417a_843c_e099_f4de_89e7_e371_b35e_ddcd;

        #200;
        key = 128'h0f7f_acb4_dac9_ffee_2954_522f_de6d_3d23;
        state = 128'h2e13_acdd_29fc_2790_7c6f_1bc3_d6f6_087f;

        #200;
        key = 128'h8683_d5aa_2ba1_4c99_98a6_6aae_3578_39c1;
        state = 128'h38bd_24fd_365e_71ad_b811_a57a_6933_1714;

        #200;
        key = 128'ha7ec_8230_bed7_bdf3_90db_2072_312b_6c70;
        state = 128'h2278_f1d6_d48a_dce4_db0a_44f9_c367_163b;

        #200;
        key = 128'hb36a_c4c2_c900_c723_778a_dd08_4fee_3f78;
        state = 128'hb333_ac7f_0a77_480f_9c29_9d43_eaa1_ee66;

        #200;
        key = 128'he047_40f6_3977_22a0_1342_372f_3bb8_0863;
        state = 128'h5f12_43f3_d66e_331b_73a8_b637_cec7_b7b6;

        #200;
        key = 128'h6969_4d73_f523_e4bd_f158_e8b0_76d9_e69c;
        state = 128'h5025_6760_b13d_a454_4116_5489_c342_8b24;

        #200;
        key = 128'h0185_1205_4dbc_163c_c1a1_cdc7_372c_24b8;
        state = 128'h516a_eb45_4783_e37a_ac63_fd03_c7b0_6df0;

        #200;
        key = 128'h0a92_146d_83dd_b006_0d61_c898_3806_80a0;
        state = 128'hd2dd_cb8a_fbdb_31f3_a85b_ed5d_f1d2_87fb;

        #200;
        key = 128'h9491_a2a4_a7cc_b94f_f947_6e13_9678_0c07;
        state = 128'h9255_2dd4_78c3_89af_c30b_533d_d419_a00f;

        #200;
        key = 128'h8011_03e9_923f_2eb4_317d_1f5b_df92_9fb5;
        state = 128'hc7af_6c0c_55ef_7753_9577_bdba_77b9_eaf4;

        #200;
        key = 128'h0047_e02e_de17_7c4c_2d40_0b7e_d237_d5e7;
        state = 128'h7f4d_76b2_2037_49f4_8d87_8858_0b52_49ca;

        #200;
        key = 128'h9fcc_c685_f009_2e2e_7494_8c44_6cc3_89fc;
        state = 128'h8e88_046b_b8cf_ade3_7ea5_428e_18f7_a25c;

        #200;
        key = 128'hc965_1f96_beb0_1b92_692b_79fc_e36c_8901;
        state = 128'h8eac_948f_a774_2f01_ee00_de7c_2e42_e9e4;

        #200;
        key = 128'h515c_c586_cb14_1fc5_6ff7_2362_7228_ece2;
        state = 128'h84e2_54b2_dc56_a031_7e9d_0ac4_40d7_cf6d;

        #200;
        key = 128'he9a1_1ea4_bd9c_0761_fd34_3c55_24b2_46fb;
        state = 128'h6b3a_ac92_b0c4_398a_b2d5_61fe_d890_e8f9;

        #200;
        key = 128'h4c6b_8444_a5be_8237_4daa_2812_0a9b_1e28;
        state = 128'h06b7_4e2f_a731_5318_0544_34d8_d827_3c18;

        #200;
        key = 128'h492a_433e_cbe4_9036_d916_3c7e_a788_445d;
        state = 128'hfbe2_9e26_274d_97f8_cc9f_ad88_c110_5061;

        #200;
        key = 128'hc947_0374_3e48_1a28_cd4d_0c6c_4d62_0da7;
        state = 128'hc625_505a_739b_4a0a_ba2c_ce60_cd5b_5fbe;

        #200;
        key = 128'h1cc1_f977_21f7_0f73_2959_300f_4ae7_6982;
        state = 128'h88cb_d7f0_23d7_ca78_1590_b2a7_53e1_0e26;

        #200;
        key = 128'h6b90_0b54_a207_639c_c850_4647_1bda_c140;
        state = 128'h6349_59ec_2966_f6ec_9e50_90ad_c2c1_026e;

        #200;
        key = 128'h5cab_081c_cf00_5c8f_9fdb_df96_a44d_128b;
        state = 128'h2fb9_2e18_3715_14d0_eca4_3245_1a46_1e6b;

        #200;
        key = 128'h18cc_d094_a267_aab2_048d_15b9_26b5_4337;
        state = 128'hf898_41f5_6361_45a8_3824_c2d8_20b8_9fbf;

        #200;
        key = 128'h08b7_9cb8_18bf_7edf_5bc1_1b13_1024_9077;
        state = 128'h49d7_7609_96e5_9c3f_6f5a_e2d7_65ea_a899;

        #200;
        key = 128'h56b7_2443_fc70_0b6b_affe_5d08_de80_4eb0;
        state = 128'h9250_1d35_f9c8_db1a_ede8_e3b1_961d_c98f;

        #200;
        key = 128'hce2c_11ac_492d_1192_dc31_7a68_bbfb_0cfd;
        state = 128'h8f04_8698_1269_38da_ecd8_65ff_c8fc_f934;

        #200;
        key = 128'h3213_3332_11e6_a72a_8f3d_47c3_a896_81b6;
        state = 128'he0d8_5163_0ed5_8a15_7b30_4028_ff96_6765;

        #200;
        key = 128'h273f_71a7_e037_111a_8cc6_0ab8_c28f_df0f;
        state = 128'h2c51_6f54_d573_868e_498c_a4c9_4bad_eb86;

        #200;
        key = 128'h9580_fc04_8121_70a8_a636_5dce_8c4f_326e;
        state = 128'h5aa8_74d0_eefb_b12f_fbcf_0e60_42e3_406f;

        #200;
        key = 128'hfd67_6287_63f2_0034_83c0_b193_090d_41d5;
        state = 128'hcdf0_2795_0335_3b3c_91d7_f83b_41ef_ebba;

        #200;
        key = 128'hb3a9_5dcf_20e1_95a8_c553_adb5_90b3_8c0c;
        state = 128'he49c_5302_fcfa_e1b5_3add_4655_8317_6ebd;

        #200;
        key = 128'h4040_cc0c_9378_a220_911c_8f10_85b1_5b8f;
        state = 128'hf8e7_a006_90f6_61d5_61d1_dc42_6115_b231;

        #200;
        key = 128'hd6dd_65bb_8eac_2bb0_c891_de53_1081_2b28;
        state = 128'hc0f6_c200_6f7e_ffd4_d3da_df44_0d29_baa9;

        #200;
        key = 128'h214e_fae4_b27b_3e76_3f4b_7b7f_5ebe_3b80;
        state = 128'h6f8a_901b_5979_9149_f5de_e135_d476_48e0;

        #200;
        key = 128'h1be6_5f72_cea1_b26e_099f_010c_5d59_d369;
        state = 128'hdd90_7192_bf0f_1ce2_0118_e24c_fecb_d224;

        #200;
        key = 128'h1506_1eeb_9fa6_08ed_d487_4be3_c48f_1708;
        state = 128'h865b_784e_fb3c_4520_7c7e_87e7_ffc9_a5c6;

        #200;
        key = 128'h02fd_e8e2_7d36_32ce_8463_c7cb_dade_8cdf;
        state = 128'h4ae4_5a1c_7066_6a43_8168_f84c_2b1b_1332;

        #200;
        key = 128'he413_8aa5_32b8_ce27_f237_3621_1789_a656;
        state = 128'he158_35e2_e249_d74f_86c5_d42a_a772_a90e;

        #200;
        key = 128'h1ce3_af0a_2e71_3f61_5a0b_c108_b800_11ba;
        state = 128'h4fab_360f_b429_8dc0_8c4d_3b45_3049_8120;

        #200;
        key = 128'hcb12_fc1a_2528_e367_5184_9cf2_5522_7441;
        state = 128'h69bf_81ff_64a9_6929_32f1_0577_cc0a_6b77;

        #200;
        key = 128'hd725_7020_0406_c7e9_82cc_f7a7_68a4_2c57;
        state = 128'hc664_7acd_0303_3c3f_6b7a_61cd_85e5_acea;

        #200;
        key = 128'h6b18_d8dc_b28a_131a_7b6c_3c0d_31de_7ceb;
        state = 128'hc29d_5873_a73d_b406_a4e5_93d1_78fe_17e3;

        #200;
        key = 128'h7410_e305_6ac9_0914_ce06_7a8a_19c1_f145;
        state = 128'h6fff_5237_36b1_1929_d61d_5a18_7784_bec7;

        #200;
        key = 128'h27dc_2a74_992f_ab84_874a_fc8b_7097_a53a;
        state = 128'hadc8_9a97_8317_a19f_5d71_9685_fcac_2cfc;

        #200;
        key = 128'hae84_773c_e4cd_7090_917f_7fe5_7a7b_ef95;
        state = 128'hefd1_2f5a_aa72_0d60_dba7_876f_88af_1305;

        #200;
        key = 128'hfc89_e0b8_1ead_81b6_d07f_6686_e4ca_a8d7;
        state = 128'h13fc_8d25_2602_f41f_5950_0711_62bb_7774;

        #200;
        key = 128'h31bc_754c_ecc0_426f_4d2a_c574_422b_85d1;
        state = 128'h39b6_6dc8_2aa4_5a8f_b555_b0f2_d8ab_0c2f;

        #200;
        key = 128'hc711_5bb5_8af1_e149_b5f0_08e7_d601_9557;
        state = 128'hc7b2_0a5c_f779_a29d_419f_0c5c_8b73_a3f6;

        #200;
        key = 128'he87e_d812_2c58_dbaa_cfd1_abf0_58bd_0b15;
        state = 128'ha7f3_9d90_dd23_0b50_eb74_9732_578a_7356;

        #200;
        key = 128'h11dd_c70a_93e4_5ee6_30c7_0ad3_7ba5_3ffc;
        state = 128'h14e4_d603_b967_1846_8f05_8516_1e11_4695;

        #200;
        key = 128'hf6b2_368d_74af_1ec3_9754_fd8b_df02_0e36;
        state = 128'h3f01_204a_ac07_b45c_5bee_e76e_7a75_0b00;

        #200;
        key = 128'hc982_1c48_edd4_5c44_664f_1894_cd1e_652b;
        state = 128'h92bf_21fa_b4be_9f1d_a54d_56b4_385b_0ad4;

        #200;
        key = 128'hf1fc_dd4c_a00b_5ed3_fa6b_7caf_5f4e_e687;
        state = 128'hc6f7_b91e_583e_5f92_3c7d_f045_c583_9beb;

        #200;
        key = 128'hc27b_7d9a_4420_f8ee_d913_ccf1_a823_550c;
        state = 128'h22de_4ebf_0491_6b41_b085_3729_0c43_16fa;

        #200;
        key = 128'h4f0c_d325_f9cc_928e_9b25_2260_6a41_608e;
        state = 128'hd297_1a93_afa4_b54b_9f74_cf57_a5f5_115b;

        #200;
        key = 128'hb0c1_c7c1_d782_ac45_85c9_d9ad_1152_882e;
        state = 128'h09ba_9486_ca45_a8d8_d567_a45d_b315_b6e1;

        #200;
        key = 128'hc266_c539_a6ef_bac0_09fb_bd19_e8c5_4e00;
        state = 128'h1127_24b3_95a5_061f_0250_f07e_f55e_1722;

        #200;
        key = 128'h9757_76e8_87fe_9e90_4d6d_0108_1236_17a4;
        state = 128'h2c1a_61b6_ae39_9dc2_26f4_0882_9ca9_f554;

        #200;
        key = 128'h082d_dada_cef1_d071_5e4c_1f26_a86b_c069;
        state = 128'h64e2_c512_3953_2525_2573_25ea_7a94_2024;

        #200;
        key = 128'h150b_aed1_7599_4118_0927_8c03_5a72_dc23;
        state = 128'hedfb_170d_b130_f1c7_ce7a_9347_199a_ad57;

        #200;
        key = 128'hc528_673e_3860_829a_4d39_4909_a251_cbb2;
        state = 128'h20ee_8213_f50a_437c_9400_ad12_300e_b34b;

        #200;
        key = 128'h77d0_332d_3230_654f_95cc_6b69_df87_6640;
        state = 128'hf089_04bf_f2bd_e520_4255_4399_675d_74cc;

        #200;
        key = 128'h7ee1_1efd_5383_94e8_9594_f9e4_47fa_d4c5;
        state = 128'hd263_61d6_1f6f_b2fd_0554_2be6_190e_ae32;

        #200;
        key = 128'hced4_b001_d42c_391e_c285_2a1f_61ae_7ed1;
        state = 128'h413a_a986_b482_e487_63f6_9e7b_dc18_a6e1;

        #200;
        key = 128'h9103_8841_9ba4_9711_451c_f9bb_15d6_4353;
        state = 128'h70e9_503f_af11_1160_646d_2a24_9bc1_ff8b;

        #200;
        key = 128'hc59b_e666_304d_b5cd_8ac3_ca64_3b5f_8cb9;
        state = 128'h72b1_db93_c452_ee37_9b63_21d6_03ec_21a0;

        #200;
        key = 128'h3cdc_439f_9afc_c894_7e06_c6a4_66fa_c1a2;
        state = 128'h9ef8_d3ac_33c6_d2a1_9ade_fcea_9a5b_b3d2;

        #200;
        key = 128'h73d2_8f08_efbe_3778_b933_7f1e_6c3f_cd43;
        state = 128'hb007_1b20_b53c_0d23_6df2_f05a_6081_43d2;

        #200;
        key = 128'h81ff_2de7_46ea_0469_4ccb_0f60_94ca_e5cd;
        state = 128'h6d3b_1fcf_4ca2_5015_106e_42e5_c90c_7cdc;

        #200;
        key = 128'h45a9_f882_01c0_6e33_0fd0_642e_3871_cda6;
        state = 128'h0d66_a162_1b88_bdb6_8dee_0c54_32b7_ccc6;

        #200;
        key = 128'h4d3c_1ee4_87ab_7fc3_bfab_4cb8_1f2b_5cff;
        state = 128'h88f0_643d_66f0_c8ad_3ec3_eee6_d9f4_cc82;

        #200;
        key = 128'hdbec_c9df_3da0_cea3_80c0_960e_c68c_14e2;
        state = 128'h145b_d95a_db8f_0f78_7d7f_4ccc_680a_04cc;

        #200;
        key = 128'h3db4_5805_4670_6925_3fc6_c792_608c_7bc8;
        state = 128'h22b5_dc36_6491_dcab_e6d7_10b3_3261_5589;

        #200;
        key = 128'h6e42_b25f_49f9_0d67_d5fc_9c5a_dda2_e175;
        state = 128'h3bb5_023f_e70f_1faa_ea38_2a57_a029_5d19;

        #200;
        key = 128'hbc8a_0ea6_a91e_7c4c_2fdb_c020_608a_6de0;
        state = 128'h5ea9_44f1_4f08_1c4b_7c27_2364_b339_5a40;

        #200;
        key = 128'hd390_6fc9_26a7_b31f_fa55_a4fb_7bdd_ed57;
        state = 128'hb61e_ff0f_278c_0843_cf53_728d_b2ce_ded0;

        #200;
        key = 128'hc45e_db23_cd3f_d8fd_8f13_6161_3aec_0957;
        state = 128'hadc7_7543_d2ba_714f_32ae_0b31_637b_8bb2;

        #200;
        key = 128'ha4c2_f7e1_3ff2_558c_c3bf_fa80_df92_ce63;
        state = 128'h7fda_f08e_c7a8_9ae8_73aa_c166_c69e_cfdc;

        #200;
        key = 128'h558f_f571_7d53_5242_bce2_08c9_269f_6be4;
        state = 128'h2e08_68f0_7308_1ea0_605e_0d3c_17c4_c534;

        #200;
        key = 128'hb653_4a8f_ea44_e26a_0df0_5997_6f30_6dda;
        state = 128'h14d6_ec37_8c3b_5243_fa2d_2560_4aa9_af99;

        #200;
        key = 128'ha3c2_ba62_c173_930c_0d60_5428_d255_3a6c;
        state = 128'h7597_c104_517d_c873_0fcc_e9e3_2f28_5b96;

        #200;
        key = 128'h24df_df3a_f709_48e5_ede1_68b7_d6d0_beef;
        state = 128'h7822_460e_73df_7521_b88e_852c_febc_c71e;

        #200;
        key = 128'h360c_1323_9267_c510_73e3_9fc1_5a58_f1fd;
        state = 128'h5dc8_a187_c878_178f_fc3d_37ae_c7b1_a2d0;

        #200;
        key = 128'h4fa3_481e_1893_a20a_6e86_1081_0321_94c2;
        state = 128'h632b_42c4_4880_fe50_2d6e_e806_c275_c492;

        #200;
        key = 128'h7d74_92a0_b0ac_156d_3e10_3511_9eed_335e;
        state = 128'h4271_4bb7_9d8b_98f8_0254_aebf_146d_a80e;

        #200;
        key = 128'h2116_662a_4390_7629_e7f1_d2d4_7824_b1d3;
        state = 128'h2210_ec7b_509d_943c_88f4_5c00_aa7d_7c2b;

        #200;
        key = 128'h51a0_be60_c592_66d9_d1f1_dece_5062_7644;
        state = 128'h5a32_e9df_f494_bf9d_aa4e_b629_c506_78f3;

        #200;
        key = 128'h18aa_b75d_da5a_8942_6c6a_275a_49d5_bdb9;
        state = 128'he03f_f02c_d5a8_ed0d_a306_ea7f_14da_84a5;

        #200;
        key = 128'h6023_fac4_acc9_afb7_5f0d_2b4a_20ad_34ea;
        state = 128'hb7ba_b087_3b41_8db2_b6ef_342c_0895_3ecd;

        #200;
        key = 128'h20ae_f694_3239_e814_ffe1_afe0_76d0_444e;
        state = 128'h55e5_aef7_0513_8709_632d_f37c_deae_5df3;

        #200;
        key = 128'h8284_c9ff_1b47_6a44_0c8c_e271_1274_1e2c;
        state = 128'h2876_aa08_3407_7bb7_9193_d7b4_5236_cde6;

        #200;
        key = 128'h027e_9310_8006_cce6_3c7d_b36b_7cc8_7238;
        state = 128'h1f52_e180_9a93_b3c0_6d7c_c209_4c78_3148;

        #200;
        key = 128'h0fda_6be6_b133_41db_4b2a_8242_6700_ed1e;
        state = 128'h144d_dcd8_dba4_203d_6ad3_b9a2_b0d0_3bb2;

        #200;
        key = 128'haa12_1f90_2d47_8aad_5cb5_4840_853c_8781;
        state = 128'h904d_ff3f_dc36_f999_755c_e797_5429_1d0f;

        #200;
        key = 128'h6dec_f415_dbdb_44b4_011a_0a9f_fb44_866c;
        state = 128'h8e3d_a483_fe45_9ec4_5b3b_2cd0_bd83_5bcb;

        #200;
        key = 128'h416e_0db5_487c_e1e7_5010_c10e_19d5_5994;
        state = 128'h0797_9277_99e3_f574_f09c_22b9_58f3_a20c;

        #200;
        key = 128'h9aa1_bd09_8f7a_8cac_8a13_470f_4e8b_97b0;
        state = 128'h7df1_0075_936a_0ae6_41f8_bb78_ff95_0ede;

        #200;
        key = 128'ha0c8_12e6_1a50_3b9f_271c_43e2_f47a_8bea;
        state = 128'heee7_0d57_73d5_9fba_319d_8ea9_0f68_2a4c;

        #200;
        key = 128'h6df4_2d3b_3d98_56ce_7bec_ceb2_dd02_8bac;
        state = 128'h8307_14f9_652e_dcf2_d7fe_91cd_923a_bd03;

        #200;
        key = 128'h1a46_911d_e941_c6f7_971e_ce4f_8185_dd87;
        state = 128'h99b6_b98d_b83f_811d_ab7f_5d1c_f2cf_02f9;

        #200;
        key = 128'h8c21_fe1b_aa2e_62f3_1001_0d80_ddb8_7580;
        state = 128'h10bd_ab54_e5d6_61a7_b5ae_79ec_921e_223f;

        #200;
        key = 128'h4f84_62ba_3999_c801_2729_ec4e_b564_23b1;
        state = 128'h4971_08a1_5757_3f77_8f2d_24b5_6cbc_534e;

        #200;
        key = 128'h3f39_4309_c0f2_dee3_a220_1dc0_c0c7_7f9e;
        state = 128'h8126_8d30_e070_e7d9_ab43_c8e7_4df4_f019;

        #200;
        key = 128'hf152_564b_7675_019c_4980_303d_bcb3_6452;
        state = 128'hc2d1_a730_ecc0_a318_8e6d_0cf3_df37_7a1e;

        #200;
        key = 128'h17a9_f6d4_6dcc_b406_5580_92e4_13b1_5d36;
        state = 128'hceb0_3bf4_77c1_8302_dadc_7286_5577_a5ac;

        #200;
        key = 128'hb37f_454f_80b0_14df_4bea_eedf_7f72_6113;
        state = 128'hab8e_4d44_8bad_e972_07e2_f229_4e0f_be91;

        #200;
        key = 128'h5e8c_e493_7aa9_53d3_f865_6c65_971c_2f88;
        state = 128'h8fe1_0b64_57ef_a136_b037_8e23_16ba_e8a5;

        #200;
        key = 128'h63f8_9b8d_e5d4_a4fe_4d99_b99b_b434_d679;
        state = 128'h186e_f973_978d_f6d8_95d1_9edc_dcca_b098;

        #200;
        key = 128'h46bd_14b7_980a_7586_f6b5_7f9a_8200_1b3f;
        state = 128'h957d_fc66_212a_1fd9_3835_2425_df8f_773e;

        #200;
        key = 128'h915e_3aa1_e0f1_3e47_c3f0_f8e6_17e7_a883;
        state = 128'h2556_3930_e1ef_19e0_6131_95a7_3991_780f;

        #200;
        key = 128'ha1b1_c4e0_1df9_3a25_cabd_495d_d0ed_81c6;
        state = 128'hd19a_43dd_ec85_53c8_f22e_f77f_5a14_3af6;

        #200;
        key = 128'h5e1c_4191_6a2b_575a_8a7a_8423_8d66_3e04;
        state = 128'h364d_59ca_b08c_963e_c632_5d85_c906_83a4;

        #200;
        key = 128'h5645_f2f5_1e1b_423d_3cf1_69f9_af65_f4d4;
        state = 128'h55f7_3b84_0431_9873_80b6_5305_5f69_101e;

        #200;
        key = 128'hd4c3_b9cd_c509_e7b0_ec20_046f_947e_8d55;
        state = 128'h8b7a_b96a_fe6d_a908_a1dd_3362_2f37_2d9f;

        #200;
        key = 128'hae3e_3c98_cea7_3ce7_44d4_9117_bf14_a323;
        state = 128'h8e8b_0293_5cab_f80c_5907_edcd_ad91_8518;

        #200;
        key = 128'h282e_85f2_f453_1a41_a63b_a8bf_ac85_39cc;
        state = 128'h4639_6d76_477f_f6fd_4a4d_3b1f_4638_3fb9;

        #200;
        key = 128'h20c4_411d_3d90_2ffc_8825_c98f_9788_fda6;
        state = 128'h9d81_422e_8c26_408c_5d48_e689_f05f_d949;

        #200;
        key = 128'h3713_b063_a4a7_b67e_9ca8_df10_aa92_d95a;
        state = 128'h841a_6055_b767_d1d0_d6ab_7dbd_5f14_b77c;

        #200;
        key = 128'h80a1_eaf5_b9ff_4967_c744_3f1a_76b0_32e4;
        state = 128'h75df_9e28_490b_c1cc_c7e0_5b5f_ffa4_3d6f;

        #200;
        key = 128'hd2e3_591b_001b_d96b_024b_e942_0cd9_e6d2;
        state = 128'hf169_103c_381a_280e_5773_dde9_2f95_d65d;

        #200;
        key = 128'h63a5_6ff7_e516_cdf4_39e1_61a3_7f4d_3545;
        state = 128'hd9b8_3907_e1cd_05b0_e5e9_df52_adba_477d;

        #200;
        key = 128'hec41_247e_e211_43fa_8905_b334_abe4_93d0;
        state = 128'h022e_e925_80e9_0ef7_331e_23a2_7f85_e5b1;

        #200;
        key = 128'hbd64_e1ae_af0a_d447_a20c_52d8_3d68_1444;
        state = 128'h1584_266f_5adc_c204_a317_c14d_d94c_00bc;

        #200;
        key = 128'h1ada_2991_be31_8d26_33ee_a3dd_5a79_79c0;
        state = 128'h3564_0461_211c_ad8e_23e5_6633_6023_787b;

        #200;
        key = 128'hd1f2_2389_0192_e199_49ca_6090_99e8_f7fe;
        state = 128'h1967_5494_c25b_8822_88f3_e059_c798_65f1;

        #200;
        key = 128'h4c0b_9d5f_76e4_f3d4_cb78_8cbe_626a_df92;
        state = 128'h9da9_5a0c_79b9_dbbe_45f8_89be_1700_a22f;

        #200;
        key = 128'h3ac7_82d2_ad86_781b_6ce1_1040_2b7e_baf0;
        state = 128'h7a46_33db_7c30_d543_b13b_55f9_24f9_1e4d;

        #200;
        key = 128'h97f8_8273_7c3d_05e4_a10b_0405_a853_11bb;
        state = 128'h140f_0d7f_523d_ceb0_d081_6d8d_17b1_d6e0;

        #200;
        key = 128'he945_92f9_919b_4e81_99b3_08e4_c94f_4d9e;
        state = 128'hbcc2_f9ea_2654_9a5b_56a5_b2e6_1372_b468;

        #200;
        key = 128'h91da_5e92_f958_1ba7_142f_b4da_3c7a_56d3;
        state = 128'h25f3_9398_a82f_3ffc_5fb5_26eb_7d02_732b;

        #200;
        key = 128'h876f_4f84_309c_ac9e_569b_3a2a_6ea3_70e2;
        state = 128'h8055_ab45_4ea8_15ce_2986_3e4a_364b_9de9;

        #200;
        key = 128'hc57e_1b95_edd7_ee26_a734_dfee_d561_5f5a;
        state = 128'hc4c6_4c73_a498_d168_1060_8650_cbab_57c6;

        #200;
        key = 128'h28cd_fd47_5368_9b1c_2cc9_f5b7_8adc_8590;
        state = 128'ha9de_6c40_7fb0_710d_f1be_b621_9ab0_124c;

        #200;
        key = 128'hdd3b_c03c_254d_5c2c_ee27_a817_61e7_494f;
        state = 128'h6235_cd3c_0e08_22ea_90af_ed20_896f_125d;

        #200;
        key = 128'had46_6476_9f83_0f52_18e3_a7a4_b001_e0c0;
        state = 128'h9703_69ae_d600_77d8_bbee_5a45_f928_0656;

        #200;
        key = 128'hf926_c2a7_acfe_3cac_4924_f1a5_6df8_b6b4;
        state = 128'h18b7_4cae_cd25_87a2_636d_4114_b975_0d34;

        #200;
        key = 128'ha447_7b1c_8e2a_8ee9_1967_3cb2_b28b_1cbf;
        state = 128'h1242_0a56_904b_0cca_8304_d0c0_ab0c_b392;

        #200;
        key = 128'hd411_19c7_c5c5_5667_d20f_907e_33b8_0654;
        state = 128'h629b_ac9c_fa3b_fa21_efa2_800f_46e7_307b;

        #200;
        key = 128'h87f5_d500_386d_14ae_68d2_ffbb_a194_b742;
        state = 128'hc01a_e13d_00bd_0ace_561a_b125_d463_c587;

        #200;
        key = 128'hd51b_2473_e986_47d5_4f6e_c9c9_b2d9_6af4;
        state = 128'h9924_e94d_b573_8597_06b6_fefb_b860_58a4;

        #200;
        key = 128'h7855_9bbd_e13b_53f8_1880_d4ac_53b3_d7f7;
        state = 128'h832f_794a_54f8_5751_5aa4_68e3_6985_7c72;

        #200;
        key = 128'ha5d4_e57a_71cb_a6c0_2b6d_6f82_acbb_dd99;
        state = 128'hc0b7_ec12_e17f_6459_4ba8_4d9e_a7db_24f9;

        #200;
        key = 128'h8d5b_6d13_68c5_2d25_ed09_73e1_ce49_57c8;
        state = 128'hb6f6_0d9c_c3aa_15c2_d755_8399_c48f_a176;

        #200;
        key = 128'he8b0_eedb_5f8a_8d12_bc35_0548_eff1_ca28;
        state = 128'h6a92_5b0d_b5fc_aaaa_c5a4_67a6_78b8_40fb;

        #200;
        key = 128'h4e3e_7f10_47a0_0145_bc4e_c389_9768_4a03;
        state = 128'h4e29_5e62_d778_4505_c046_2c8f_35df_47a5;

        #200;
        key = 128'ha56e_73ba_f1f8_3395_c720_d5a1_bc88_b1b6;
        state = 128'h5859_0d0e_7590_5601_31a6_1edd_ce0e_62b6;

        #200;
        key = 128'h68a1_0334_849c_8703_2819_0777_eebe_77cd;
        state = 128'hda4a_44b8_824e_63ee_021e_127d_08f4_9a9b;

        #200;
        key = 128'h4365_b7dc_21ca_82b2_5879_a57a_9178_ea6a;
        state = 128'h8d74_ed90_4b9a_9468_03a1_db4a_7439_5311;

        #200;
        key = 128'h8d9a_3744_a6fb_cd62_ede1_3cdd_fc8f_7c9b;
        state = 128'h7dce_bbcc_e931_09c9_edc5_ca21_3d26_bf92;

        #200;
        key = 128'h6d76_6fb9_d743_996d_7f35_9843_1eaf_e8ac;
        state = 128'hd557_ea5d_67de_a501_7afe_b637_d5f6_4bb9;

        #200;
        key = 128'h6a78_3a27_2a22_3813_97ea_7916_74df_95c0;
        state = 128'h05f2_8a74_d588_a96a_a90e_9703_1991_cb8a;

        #200;
        key = 128'h76cc_a152_4860_3078_049b_1e87_bc5d_9240;
        state = 128'hecb9_c074_7c6d_5af1_023d_4087_7c90_9c85;

        #200;
        key = 128'hb870_44f2_b07e_1acb_d83b_78d9_4103_4e1e;
        state = 128'h9f82_b933_bc07_076a_b6a6_d19e_c452_ebc4;

        #200;
        key = 128'h3a15_0d31_41c5_554a_0003_ef9d_829b_c009;
        state = 128'h29b2_5124_f017_0955_52d9_29ba_0c69_e904;

        #200;
        key = 128'hf543_a47c_4455_2317_d8c6_7213_a338_87a7;
        state = 128'h7b14_c713_4364_d0d6_1dc4_01fe_4a34_c957;

        #200;
        key = 128'h0728_f667_5a87_0b12_4132_5085_7044_0adf;
        state = 128'he202_950d_36de_dabb_8741_5cea_f98c_877a;

        #200;
        key = 128'he8ab_6839_0869_5d4d_226d_e94f_d49c_e05c;
        state = 128'h094d_e5d5_2b21_6fbd_9c2d_4ff9_5ae1_bb05;

        #200;
        key = 128'haeaa_b68e_afb3_5902_f86f_74b3_1414_35aa;
        state = 128'hea77_345a_5a91_aa9b_c295_ea29_61b2_5d70;

        #200;
        key = 128'h9f8e_437f_7fa3_d7da_922c_8da4_7be9_2e96;
        state = 128'hcb2a_0fef_edbb_49f2_90dc_7cf4_f805_f2b5;

        #200;
        key = 128'hf053_7760_e5ed_84d1_8899_7771_8c70_ee75;
        state = 128'hd632_8eea_cec8_d74b_289f_09ef_6e54_4038;

        #200;
        key = 128'h468e_bd5e_5bbb_eb74_204c_de15_81c5_47bb;
        state = 128'he2ed_74be_8b41_5e5a_e4b7_827b_83a8_2bcd;

        #200;
        key = 128'h5f2c_fd1f_a629_94af_067d_2bb7_2734_4872;
        state = 128'h226a_62d7_a1c7_4af1_2844_1f5a_386b_ff6f;

        #200;
        key = 128'h1b11_79e2_9feb_8763_f332_a7ce_15dc_6246;
        state = 128'h02a3_e451_e471_4827_4c23_495f_0ebe_c91f;

        #200;
        key = 128'hd2c0_5f88_dfe0_30a5_4720_c0c6_72be_8eed;
        state = 128'h79c7_ac77_58c9_2bf1_74ce_9245_c08a_d082;

        #200;
        key = 128'hf94d_bc88_ec2a_7991_be73_400a_8414_ced7;
        state = 128'hbf9a_602c_31a0_b9c7_50b6_9b23_b499_5db2;

        #200;
        key = 128'h6168_1a51_1d0d_1f93_81ed_adb4_e438_93bf;
        state = 128'hefed_38c3_9360_76aa_14c4_2d52_597e_c39f;

        #200;
        key = 128'h4096_5d69_2ac2_6e5c_8682_39ed_54d4_7a35;
        state = 128'h3d0e_2707_2bfd_f36b_24bb_3e81_951b_d25a;

        #200;
        key = 128'h35b8_ab44_4452_5cf9_f8c2_b286_d291_c3f2;
        state = 128'h08ce_62c8_0027_2cae_9a88_f85f_05fc_8ee1;

        #200;
        key = 128'h1f6e_4fb4_0f28_e7e4_6f9a_d369_fd73_38e8;
        state = 128'h9ce0_c232_4935_f162_9992_a382_79f9_2b3c;

        #200;
        key = 128'h19de_f202_159a_17e6_dfa9_1499_f166_a508;
        state = 128'hd892_252d_3a1e_02a2_aa67_5671_2519_716d;

        #200;
        key = 128'h59d4_7e42_aabe_a1dc_ac5c_e3d8_b5a8_6400;
        state = 128'h5b30_3818_8f0c_3577_9a5b_9f7a_ece1_d4f1;

        #200;
        key = 128'h13e2_d235_cb65_ddc6_e901_197d_8689_f911;
        state = 128'h148b_7649_4e8d_b083_67c1_7081_058a_ba96;

        #200;
        key = 128'h6e68_dbb8_8e51_a28b_ee39_59ed_4922_4e6e;
        state = 128'h7538_e08e_5283_c8ec_67c7_10bf_0093_d2fe;

        #200;
        key = 128'h323c_be5b_2801_449b_4951_28db_23ef_2891;
        state = 128'h4e8a_c997_93e0_4cdb_ef19_aa93_9247_e116;

        #200;
        key = 128'h1278_c416_b821_1f27_c731_4e64_0139_1f02;
        state = 128'h65ab_79c1_4b13_e805_dcc1_dfd4_5e01_e88e;

        #200;
        key = 128'h73f3_33b0_390d_8ba3_20aa_d39c_7f5c_21a5;
        state = 128'h4eab_10db_27ed_4fa9_5b61_6a99_6309_af9b;

        #200;
        key = 128'ha8f7_91b5_53fe_9176_dffb_2414_5c77_c9d9;
        state = 128'h5b26_8ea8_9047_0d0e_5a06_cd80_0a2c_b0e2;

        #200;
        key = 128'hc550_5132_13bb_e356_1f76_75a2_d023_2fb4;
        state = 128'hb278_6249_687e_7c97_f231_fcd4_4b23_ccad;

        #200;
        key = 128'h6c46_2d0d_c523_b12c_98c2_6c6b_b878_3e3e;
        state = 128'h50b8_8a8b_50b1_97ea_e611_2217_0acf_a499;

        #200;
        key = 128'h1ebe_9d1d_5bdc_b614_f21d_1a7b_049c_3514;
        state = 128'hcdb4_5914_b710_51bb_5969_2cbd_2c12_79f3;

        #200;
        key = 128'h298a_dce7_7b95_f381_a82a_72b3_76ac_13d9;
        state = 128'hccc9_201b_9764_a32d_1577_65e2_262a_e41c;

        #200;
        key = 128'h227f_298e_e68e_3321_0128_aa1d_f799_1ea6;
        state = 128'h2f1b_d4f7_c2f4_9835_585e_c81d_068a_b375;

        #200;
        key = 128'hbe41_b862_9f83_9245_c1c3_4f20_e362_ba62;
        state = 128'hb660_4e3f_a24e_dc14_630f_b58d_7f4a_9474;

        #200;
        key = 128'h7a79_5a7a_3868_e473_3e9c_0250_cf06_d8a4;
        state = 128'h0013_e2f6_da19_481c_e211_39b1_fe91_12cd;

        #200;
        key = 128'ha79b_753f_4254_a23f_6007_2a47_0706_4752;
        state = 128'h32e8_8b83_3365_96ab_10b5_58d8_ea6d_1c8f;

        #200;
        key = 128'h2779_9863_921b_b6a6_4b34_bf24_4ab9_66f4;
        state = 128'h2213_9dcb_9057_a5a6_48cf_5df8_f31e_f6a1;

        #200;
        key = 128'hd606_2917_877c_40a5_153f_574b_2400_107d;
        state = 128'h021a_7c5e_04ca_3429_90bd_087a_bf36_fd7b;

        #200;
        key = 128'hcd20_f315_d32b_9988_34f5_b586_f775_c6c8;
        state = 128'hed7b_b126_43c9_c21e_74f0_a35e_a87f_1335;

        #200;
        key = 128'hda37_1f88_379c_4032_e10d_b84a_7d64_9af6;
        state = 128'h48a7_42cf_416f_565d_7d1d_dcdb_d264_00fb;

        #200;
        key = 128'he95b_b47e_536a_4242_19d2_d928_a06e_ae92;
        state = 128'h8583_9139_5cd4_8390_c741_fdc0_81ae_c028;

        #200;
        key = 128'h61e7_955b_7156_9097_a439_e845_a4ff_e714;
        state = 128'h5cb1_e023_274f_b222_84a3_a78d_40ac_6003;

        #200;
        key = 128'hdd57_d21e_9ceb_ee82_5ded_d8e3_8321_b3fe;
        state = 128'h57fe_925d_b545_2294_d991_18a0_d58e_9cef;

        #200;
        key = 128'hefff_a504_8e01_dd4f_2732_48d8_f3f5_acb3;
        state = 128'h76ce_4980_7d4e_3002_2bb3_7c46_c479_0d56;

        #200;
        key = 128'hc8ba_76e6_afcf_1aaa_70d1_7309_e423_3ef8;
        state = 128'h272b_dcbb_e2cd_ee46_352c_2693_8ed4_b6c5;

        #200;
        key = 128'hd2bf_539f_36ec_a5f5_24a0_6b54_0ae0_8fdb;
        state = 128'hc7f0_6c8f_d2bf_30cb_ca21_3104_640b_9313;

        #200;
        key = 128'h3ae7_6b3d_773e_e641_fde6_b85d_2154_f9f7;
        state = 128'h2757_5fea_c353_ebd3_a847_e5d2_bbe8_9e7a;

        #200;
        key = 128'hdfa0_6fd9_4f10_909e_4616_10b0_6e67_4951;
        state = 128'h6c90_0df4_3720_7799_b774_21f0_29db_8219;

        #200;
        key = 128'h9f1e_5b2b_492c_0acb_f3ed_cd0f_000c_321c;
        state = 128'h5e0c_55a9_b684_8899_86db_c87a_192d_bfdf;

        #200;
        key = 128'hc6e8_715e_32b2_c704_c525_e635_7072_d6be;
        state = 128'h0055_5458_2ec8_c54b_fd97_23fa_5599_22ad;

        #200;
        key = 128'hdc21_bfbb_535f_397c_5e6d_0373_95db_9c5e;
        state = 128'hdd97_1fee_28f2_dfdf_cf43_5104_3be3_4ea2;

        #200;
        key = 128'ha424_bc45_d14a_9eb8_4c90_1d06_3c1a_493b;
        state = 128'hd46e_53b2_1f33_4599_5ea6_04bf_c5a4_56c4;

        #200;
        key = 128'h27ef_7c99_a60c_58d7_096a_09ca_3a32_ea33;
        state = 128'h022d_1434_346d_5e2c_66be_6f96_0f47_0e62;

        #200;
        key = 128'h7b64_a0e1_8a21_83c4_62f2_46fc_d09b_fc6f;
        state = 128'hd3aa_a60d_417b_32c4_152f_d978_2af9_e259;

        #200;
        key = 128'h9f11_ebe0_749a_69cd_b508_6fee_8824_bbd6;
        state = 128'h245c_53da_6a21_f5e2_29bf_19d3_d4bb_428a;

        #200;
        key = 128'ha3ca_2171_f4c1_d494_1da0_f428_a007_7203;
        state = 128'h9673_d30a_d886_f85e_9468_023c_9ecd_c5fb;

        #200;
        key = 128'ha11c_3c91_ac0c_d550_a94a_96a9_0d46_91ac;
        state = 128'h0fa0_661e_d877_edee_71eb_ee65_ef53_59d3;

        #200;
        key = 128'h62a8_36d6_0c39_4e17_effa_5bc5_4601_1c0a;
        state = 128'h2d4e_1f8a_6900_d643_d296_73fd_6b48_738b;

        #200;
        key = 128'h4110_9389_3ad5_0181_662e_d9d5_af9f_f0b6;
        state = 128'h4c56_59ec_81ad_2928_647d_3da5_3a4a_e5e2;

        #200;
        key = 128'ha99f_78aa_6257_d543_0085_b593_7478_22f9;
        state = 128'he65e_9bd2_2b65_413e_8119_e5ce_adc4_162e;

        #200;
        key = 128'h10a8_af6f_413e_ae07_8f63_d647_c16a_b07b;
        state = 128'h486c_3546_2034_9ef5_ff81_8f2c_2be9_ea0f;

        #200;
        key = 128'h82d3_4606_d0d1_c694_1f50_b699_6ac9_d585;
        state = 128'hf6ae_8299_ce1a_0c1c_b77c_755a_97db_fa92;

        #200;
        key = 128'h9499_0ed5_dcdd_3477_925b_eaa4_c37e_33de;
        state = 128'hac24_c141_38bc_7232_bac2_ad3d_def4_ed05;

        #200;
        key = 128'h3cac_3757_f5cb_80f9_151f_5cff_9c40_5e10;
        state = 128'h2ebc_caec_a7be_6bb9_7321_4ce7_4575_65c7;

        #200;
        key = 128'hab88_16c9_7574_4757_0851_3b12_d14b_0d30;
        state = 128'heb93_4ea8_75ba_d7bc_2418_500e_7404_1922;

        #200;
        key = 128'h94e2_30ca_09e6_2693_c2a5_d32b_2880_7094;
        state = 128'hc059_6267_1f4b_0143_11e8_a524_fac2_980f;

        #200;
        key = 128'h5c51_b5ff_e48a_9188_45bd_d6f8_b3bf_1ccd;
        state = 128'h6c00_bb9d_a73d_2c81_61d7_0abc_6219_34d6;

        #200;
        key = 128'h4238_82e9_e042_c65d_3f08_520e_1324_a6dc;
        state = 128'ha829_2a27_8977_aae9_cbbc_0dc4_67de_e7a8;

        #200;
        key = 128'h3013_e416_5412_b7a2_09dd_a23f_1eed_28c1;
        state = 128'h46b4_1ac6_d544_4ce2_024a_ec70_db28_0ab0;

        #200;
        key = 128'hb5d1_0426_806a_faa0_f6ac_c969_3911_faa2;
        state = 128'h2c6b_dea5_4eb4_51f0_73b2_2b8a_74ce_b656;

        #200;
        key = 128'h8ee3_9a7e_5e26_e7b8_58ba_209a_ee68_af5f;
        state = 128'h5d01_6377_ca09_805e_de10_9337_5327_8672;

        #200;
        key = 128'hcd83_0de3_a8c4_ba81_38f1_a0bc_b5ce_1e3d;
        state = 128'haae1_df4b_e1a0_4008_1123_8831_6586_155c;

        #200;
        key = 128'h31ff_fb2f_b3d5_5311_66c7_0f67_1929_ace5;
        state = 128'hc539_39be_8fe3_3237_dc22_3751_33c7_99b1;

        #200;
        key = 128'ha2ca_07ee_fbfc_37d1_e141_c2ab_d37e_2c2d;
        state = 128'h87ca_c1c5_3479_851c_3d09_31ae_0efd_eca0;

        #200;
        key = 128'h0b35_51ab_cdbb_aa01_47f8_c848_dfc8_ca47;
        state = 128'hfcf9_804e_3562_f5c0_c00a_e498_4725_b0e8;

        #200;
        key = 128'h1fb3_9642_9326_947e_422f_4ea5_a9bc_fe4e;
        state = 128'h5f57_3aec_3f97_54e0_d883_f94f_0cd5_f7ae;

        #200;
        key = 128'h3447_35b7_0e0a_c97e_8514_cd98_edfe_cf1d;
        state = 128'h2408_fbd2_5051_6367_fb2e_b4dc_cda0_a3c9;

        #200;
        key = 128'haa92_b3c6_c6f9_8bca_fbb2_8248_b043_b458;
        state = 128'hd5d5_7210_4144_8bb1_4136_c220_a6fd_af7e;

        #200;
        key = 128'he112_a8b1_e8e0_f866_23cb_87f8_7de5_3614;
        state = 128'h6eb6_bd35_d28c_211b_a986_f95e_fd92_9a57;

        #200;
        key = 128'hd780_dd8a_1a81_ee51_343a_9069_b908_d5c5;
        state = 128'hd908_556b_5b33_0bf3_0d28_439a_8806_2c83;

        #200;
        key = 128'h5ce4_ce06_c9e8_1228_3852_ea95_b09f_1ea6;
        state = 128'hd69c_62b5_c3d9_3d6c_c071_8132_4c3c_cab9;

        #200;
        key = 128'he34c_0320_e2b3_44b9_1d9a_9dba_016e_3a2f;
        state = 128'h0526_659f_bd5d_2d2c_62cf_5922_23a5_b38c;

        #200;
        key = 128'h30bb_d41d_5163_cc40_ead0_7074_afba_5ba0;
        state = 128'hd5c9_2cd4_daf3_76e0_fccc_fb06_6388_9b0e;

        #200;
        key = 128'h6bcf_3090_a0d7_4b88_7274_99f4_3216_5b42;
        state = 128'h4e94_314c_8374_6fc6_eec0_bee0_4ae3_cbf7;

        #200;
        key = 128'hbfd6_e7dc_d7d3_1ff1_13cf_46a6_4d13_c54c;
        state = 128'h43ec_82be_979f_9d68_4a4e_400b_f6ec_9545;

        #200;
        key = 128'hdb50_c5ef_cfdc_a8ae_b0a1_aee7_afe7_ec50;
        state = 128'h3556_1aa6_02df_deb0_74f4_2082_ba09_bc31;

        #200;
        key = 128'h828b_16f1_ae04_097d_e88e_2f7c_f63d_a5ea;
        state = 128'h5f32_58e8_96cd_3aad_0f91_f218_d7b5_2188;

        #200;
        key = 128'hb816_a42e_4ab9_47ee_a22c_24cc_0aa4_abcc;
        state = 128'hcb88_0272_8605_ca4c_475c_7088_5482_21b2;

        #200;
        key = 128'hea01_08de_27e0_0174_dfbc_f9a4_c085_9ce9;
        state = 128'hafdc_86b5_fbe0_03ff_50bb_1b56_dee4_43b6;

        #200;
        key = 128'h5506_4718_21d4_d884_d06c_c35b_9eea_a6ad;
        state = 128'h1ab0_1ba4_090d_5d3e_d789_9a43_8809_97a0;

        #200;
        key = 128'hfb78_583b_114d_3584_0de8_2432_9537_647f;
        state = 128'h4665_1df8_1fae_1fef_3198_edb9_8ab0_beeb;

        #200;
        key = 128'h4fef_ea43_f01b_cba5_51eb_fea3_65f8_f227;
        state = 128'h8911_1953_62fa_d5fa_b463_8d10_95b5_af8c;

        #200;
        key = 128'hffea_d455_8d4c_ccae_3f5d_5d6e_e59d_856a;
        state = 128'h4e3e_d0a8_7aca_68bc_ed34_0154_99e8_a723;

        #200;
        key = 128'h48ed_3f35_2dc9_5599_98c6_6ae5_d9fd_228a;
        state = 128'h946c_6ef3_c824_558c_1833_9d3b_14c1_56a7;

        #200;
        key = 128'hdf7b_f3a4_9d6c_4ef5_ffec_d57a_27dc_46ad;
        state = 128'hfda1_dc8c_9abf_f192_17af_d61e_4fa5_da86;

        #200;
        key = 128'h83e3_dc43_6e71_dbef_3a15_cb3f_085e_299b;
        state = 128'hcb0b_92f3_2d81_5806_3cc7_516e_a4d5_1dcf;

        #200;
        key = 128'h4395_8209_734a_4fc9_42cf_ef15_0f01_c6e8;
        state = 128'h5d8c_78d8_8c07_bbad_066d_3f8c_7039_61fe;

        #200;
        key = 128'hdfa6_34f2_59fb_a8e1_a548_3312_46a2_749c;
        state = 128'h3bdd_f495_12cf_5e0f_b637_b82b_6401_84c4;

        #200;
        key = 128'h6e8b_aaa0_7e92_dd5a_9c58_a001_62cd_c17b;
        state = 128'h03da_736b_fead_3757_10b5_1f66_5d2a_212d;

        #200;
        key = 128'h1999_2697_bc3e_c974_a4c7_4ac2_1193_c66c;
        state = 128'hd121_9129_004c_2345_ed6e_3df2_49a3_83a8;

        #200;
        key = 128'hf1a6_4173_101b_f5da_fff2_0b1a_92bd_d114;
        state = 128'h2530_205a_77af_86c9_55fb_99fa_81d3_dbae;

        #200;
        key = 128'h3d24_141f_3e4e_7d39_f618_6be2_0049_1c65;
        state = 128'hc704_a661_7733_e2fb_0663_a047_5868_8e53;

        #200;
        key = 128'h2a0e_8e6f_69dc_1fc6_9404_2a5f_39ae_0cd1;
        state = 128'hc4c0_6404_6809_c8cb_4c9b_3259_6f7f_51fc;

        #200;
        key = 128'h0d38_a6f5_3059_d985_9f2a_80aa_cc32_475e;
        state = 128'h5c2a_b566_6ba3_4b3f_1635_db01_f51e_6db2;

        #200;
        key = 128'hb91f_c0db_973c_7db6_0d61_daa5_6c50_a4a5;
        state = 128'hb41f_ee03_37b7_ddea_04ed_ddd8_2985_45bb;

        #200;
        key = 128'h0365_f7cc_0d0c_0b37_b242_6e5d_7508_f936;
        state = 128'h6d39_5e5d_38b1_12a7_e76f_20b4_c5c9_57f6;

        #200;
        key = 128'h86b7_086b_ea50_29b1_3b5c_f768_8d28_aa84;
        state = 128'h0caf_adb6_8394_a452_3f37_4b45_b56f_d14a;

        #200;
        key = 128'hced0_8a42_c31d_da69_8d1a_f09e_40a5_4892;
        state = 128'h9b0a_a262_f329_91d5_4486_96e4_fce8_ca90;

        #200;
        key = 128'h7b70_03e0_b78c_99f3_2599_2a10_579e_64ac;
        state = 128'h05e1_e3c7_08de_205e_ad5c_4add_68c7_17b3;

        #200;
        key = 128'hdd11_f15b_a4d4_84cd_a9e6_34be_7a41_740b;
        state = 128'h899b_4401_92bf_8ba6_3ffc_f643_5f4b_aebc;

        #200;
        key = 128'h1db4_b8e8_cd38_9c39_860f_9f55_1a1e_367a;
        state = 128'he7a6_e0ea_21c1_5402_95d2_3c1d_112b_2522;

        #200;
        key = 128'h77e9_7a26_649d_af31_636c_99a8_66a6_350c;
        state = 128'h0960_fb0e_5aee_ea10_a180_1e37_2228_77db;

        #200;
        key = 128'h981b_1632_40ff_61d5_b621_ebc8_9f64_0a1c;
        state = 128'h96ce_e916_8998_4a57_c086_09e4_be11_cf6c;

        #200;
        key = 128'h3ffa_5975_d4e7_bbba_1b62_607a_663c_3d3f;
        state = 128'h272a_2df9_9f70_cf31_2103_d4d6_5ccb_3a38;

        #200;
        key = 128'h036c_b671_63b0_cb4e_9e97_348e_a661_1b09;
        state = 128'h189c_7476_0238_f987_3b01_861c_6167_931e;

        #200;
        key = 128'he627_c8b1_eadc_cb2e_2295_3eef_c98e_0a2a;
        state = 128'h04b2_fc16_e131_15d1_587e_0c9d_7b81_b794;

        #200;
        key = 128'h8100_e621_5482_3aa8_ed4a_196a_829d_ef7a;
        state = 128'h6be0_2c87_effb_8adf_2179_c78e_03fe_4ab6;

        #200;
        key = 128'hbc78_f700_1425_9ffc_9661_aa9e_9ff7_1759;
        state = 128'h244f_b9c9_0e09_1882_468c_93b8_ebbf_ae75;

        #200;
        key = 128'hcc97_c027_371a_515b_d519_5e98_34b9_07c8;
        state = 128'h8b49_d84b_2bb3_2b4c_c088_e41e_8ca2_3804;

        #200;
        key = 128'hc0bb_c864_1cb9_3758_c801_208a_9372_52c2;
        state = 128'hf0e2_d60e_c2d8_2364_2b11_4f23_c333_358b;

        #200;
        key = 128'hf461_c0b9_d3c7_1baa_9230_9bba_28b4_1369;
        state = 128'h6b17_5a58_3689_591e_5fe4_1041_1dce_6c77;

        #200;
        key = 128'h2041_9d33_8397_94f6_3ed5_8064_80f1_7327;
        state = 128'hc754_153e_022b_d8e1_7d0f_c494_af67_3bb0;

        #200;
        key = 128'h3ffe_7f8a_ff48_99c3_fa4c_392e_2a0e_4df5;
        state = 128'h154f_42d7_08d9_a2e4_c8e9_fb6c_a3c1_1d45;

        #200;
        key = 128'h0656_f651_47ba_d5c2_8824_dcdf_48cf_64f3;
        state = 128'h8143_38f7_1173_cc0b_81c3_6eff_318d_c1c1;

        #200;
        key = 128'h1a6e_a86a_3cfd_1575_c52d_94ef_9d18_1316;
        state = 128'h6264_a849_9501_a937_de09_0982_e290_0dd3;

        #200;
        key = 128'hf6cb_97c0_dd48_7ecb_929b_3538_e073_893c;
        state = 128'h6934_cf09_d930_ad6f_8598_e7d1_4abd_cef1;

        #200;
        key = 128'hd6e5_f05d_541b_b024_a542_2437_8465_58c3;
        state = 128'hf4e6_347f_a46d_f616_bdcd_6e82_5b39_e1f8;

        #200;
        key = 128'h7efd_d0a5_5982_159d_b5f1_ac7e_aef9_0404;
        state = 128'hf729_f3bc_acc0_647b_2b0f_3a05_787e_46b1;

        #200;
        key = 128'hf572_dbd0_5867_f77d_4b67_a930_261b_4713;
        state = 128'h5221_bace_2cbe_16be_5391_0bdf_de50_f828;

        #200;
        key = 128'h9a1d_ba55_efd4_6242_11c4_50ea_ab88_38d8;
        state = 128'h76ce_7c81_53f1_345e_3491_40a7_7600_87c8;

        #200;
        key = 128'h9ef8_0ffc_7e38_8a95_f213_2a40_a119_87f2;
        state = 128'ha57d_e062_348d_6d92_9480_093e_3c53_0493;

        #200;
        key = 128'hc497_0287_5481_4645_8277_df84_8582_43c5;
        state = 128'h6296_1b88_dbd1_3aca_acc6_00c7_a7ee_3b08;

        #200;
        key = 128'haed0_6b7f_7679_a96b_4cdb_f047_f7c2_b31c;
        state = 128'h40b3_c405_52a1_6f96_5867_80a0_ae1e_d59f;

        #200;
        key = 128'h0226_90af_8cf9_b789_0ea8_47db_9c10_4b9c;
        state = 128'h9236_025a_a1c0_df15_ca89_fa2e_0bdb_f70a;

        #200;
        key = 128'h679d_b7cc_5272_c3f3_5d2d_f300_7736_f920;
        state = 128'he4ab_3f8a_83c5_0f2c_31c3_3140_d1d6_5ebf;

        #200;
        key = 128'ha7d1_de36_9bef_596b_2dc0_e6ae_c69d_96df;
        state = 128'h2f2d_795d_7a38_a298_bf29_45bc_1148_560a;

        #200;
        key = 128'hd38c_efc7_3fb7_8bac_7add_7d12_f3bc_3b27;
        state = 128'h11c6_6ac1_c0f0_a415_deed_114d_8aa5_0d52;

        #200;
        key = 128'hdec6_211d_5102_d4f8_2ab5_14cd_67f2_fa40;
        state = 128'h462a_6104_c078_75b7_82cb_d8f4_79f5_10c8;

        #200;
        key = 128'h1ce6_f248_839b_1b02_1ad2_0aaf_86bc_67b2;
        state = 128'he62f_75bd_df7b_2daf_9ccc_0553_ea56_acea;

        #200;
        key = 128'h4c91_aa34_381d_95e6_3bc6_ffa2_714a_270d;
        state = 128'h8d0e_20c0_fb81_7172_0764_8928_4f31_d7bd;

        #200;
        key = 128'he2ea_baf3_88ae_f59e_a6cc_d676_dccb_f1f9;
        state = 128'hd18b_6e9d_8c8e_e968_c570_7a82_8aed_a511;

        #200;
        key = 128'hca8a_4253_30b1_b0ba_5ef1_828c_7a62_6ae7;
        state = 128'h03a4_0ba9_9f6f_f549_2132_820b_6d56_ee8a;

        #200;
        key = 128'h9540_d4ea_7f80_1ddb_922d_db6c_114a_e6b0;
        state = 128'h87c4_9e16_8712_4cd7_8fa1_3c4d_97c8_b89a;

        #200;
        key = 128'h43f7_71a3_ac76_8c81_9589_c0c5_6d33_bfd4;
        state = 128'h783d_22b4_9eff_f5ab_5895_abb5_d4bc_07a2;

        #200;
        key = 128'hc78c_80a1_ae5c_9457_da2d_60dd_5572_5ef6;
        state = 128'h6f22_9fad_a8c4_efb2_09bb_6b22_20db_f0c6;

        #200;
        key = 128'h28ff_398e_41df_9f64_26cd_cc0f_4697_186c;
        state = 128'hc898_9cd8_c978_3e1e_45ce_385d_8116_38de;

        #200;
        key = 128'h9eb8_4d99_80d7_8e23_0f42_c356_19fb_eabc;
        state = 128'hf2ee_37cf_4b58_cdfb_fac8_9147_81fb_177f;

        #200;
        key = 128'h2545_aa34_4e21_8ecc_8a2d_1571_6f51_0256;
        state = 128'hf8f7_9298_ba8f_287a_e97f_ab44_a078_d719;

        #200;
        key = 128'h8e93_4d80_36b5_2900_483f_fdc9_8b49_5e1b;
        state = 128'h733b_c559_7aa2_8187_32a2_32c9_aab4_ff29;

        #200;
        key = 128'h382d_bb6b_c24f_e79c_1a1b_cbab_bcbc_4b5f;
        state = 128'hf89c_5947_ff4c_06c7_9bdd_f539_6d71_20b6;

        #200;
        key = 128'hce5f_da02_500b_7096_ebcd_828e_01ae_01a4;
        state = 128'h640e_82b4_b85e_010e_6a0c_0351_0112_d45d;

        #200;
        key = 128'haeb4_a45e_dd71_101b_66b2_3fd8_b70c_8779;
        state = 128'h971d_d32f_5408_5f41_11b3_c6b9_fdc2_3f26;

        #200;
        key = 128'h1afe_5081_79f1_49a0_f24e_8ca6_6a45_0563;
        state = 128'he91b_2193_aee7_1e09_1c95_f5b6_d93d_3aec;

        #200;
        key = 128'hf483_12c3_48f0_5932_839b_3965_e786_62fc;
        state = 128'h77ec_587b_d7fd_f20a_b590_0ce8_cf34_37cf;

        #200;
        key = 128'h1ac7_3600_65eb_99bf_70a9_0e28_8e3e_b72c;
        state = 128'h2e70_c7c7_296a_4304_516c_88d1_2607_4ae0;

        #200;
        key = 128'hd9b4_47b1_9e56_9069_353b_c5a8_0344_0015;
        state = 128'h48fe_52a3_7dd3_1106_fea0_8f59_a79c_80d5;

        #200;
        key = 128'h5365_7ba1_37fc_db9f_7d24_9427_d243_b4ff;
        state = 128'h7c2e_ba1e_bd79_7def_d2f0_1c60_319b_55a6;

        #200;
        key = 128'hecaf_533d_6865_e038_1a98_32ae_13c5_33c5;
        state = 128'hefec_b60d_c3d1_bb96_05d6_a0f1_cb8c_c4d2;

        #200;
        key = 128'hdf9a_3e39_4b04_5f72_b7e7_62fe_45f4_ecc6;
        state = 128'ha7fc_bd9c_55fd_da7e_a1aa_bbc3_cc44_6372;

        #200;
        key = 128'h702c_659a_f686_4edb_e445_c37d_4d42_5ad7;
        state = 128'haac2_7924_f4f9_1057_176b_69ce_06df_37e4;

        #200;
        key = 128'h4596_5aca_5903_2e3d_82c2_d51c_0aee_265e;
        state = 128'ha254_3dd7_1c66_be4c_94a2_9062_b07f_0da3;

        #200;
        key = 128'h4f00_6b45_3d5d_e55b_8198_56b7_768b_4ddc;
        state = 128'h5455_ec7b_354e_bc61_82d2_564a_7c1d_4493;

        #200;
        key = 128'hf6ac_0af8_6e23_6504_45ab_de22_4d8a_fd2e;
        state = 128'h9127_eb9c_bb98_bb7f_743a_9b1e_1145_2095;

        #200;
        key = 128'h0468_fdb2_cc06_fb44_3ec9_4b1d_f374_9994;
        state = 128'h0f55_8c0a_e5ea_4e8b_fdc1_3d20_0f7f_3640;

        #200;
        key = 128'h7c74_a586_8c70_0e17_2c8f_a2e8_22dd_b342;
        state = 128'h558e_2ff2_a73c_7484_b103_6511_a733_9f90;

        #200;
        key = 128'hf452_c329_f125_36b1_4d70_404a_61fd_496a;
        state = 128'h5bac_6c37_0712_68a1_1ef2_ad8e_94d2_b934;

        #200;
        key = 128'h98f2_1331_dcea_d3bf_7e7a_e248_1316_db90;
        state = 128'h1c09_e719_3ef5_25be_7140_711e_8d43_35ff;

        #200;
        key = 128'h8807_e00a_b873_2281_4ae0_bfda_75df_fa24;
        state = 128'h6723_e38b_a0e8_14e9_a7bf_326b_69d7_cdad;

        #200;
        key = 128'h90c9_184b_8dbb_07ed_53d3_b67e_0498_2099;
        state = 128'hc8b4_696d_4b48_d32a_c6c9_7fab_8571_7a44;

        #200;
        key = 128'h0570_ccd8_aded_b348_554e_f3d4_1b2e_2097;
        state = 128'hd98d_8722_8cba_77ec_de9e_4204_f3cb_00c7;

        #200;
        key = 128'h6339_4ec2_c5cd_35aa_972e_c2df_8139_a354;
        state = 128'hc815_485f_4867_a508_ea3e_7914_d406_e7eb;

        #200;
        key = 128'ha123_0e38_152f_9006_f50e_918d_63e3_f5a5;
        state = 128'hd2d1_8f64_83b0_bc61_b2b5_943f_2159_2dc7;

        #200;
        key = 128'hd163_0ba3_580e_40b6_6091_0349_add7_786e;
        state = 128'h42e5_3bc8_4e93_2ef6_8afa_6bb4_9fb6_ca25;

        #200;
        key = 128'h9d9a_423a_7a06_fe79_48e8_80a4_88d9_cc60;
        state = 128'h5235_707d_9d10_e1ab_763b_58f7_b586_fb4c;

        #200;
        key = 128'h0fff_a612_cd3c_c7bd_ed50_eb03_c2f3_65a7;
        state = 128'h0cb5_b2b2_aed8_2e9e_d53b_249d_2616_0cc1;

        #200;
        key = 128'h9f6b_626f_3b48_a597_7306_a720_3064_f310;
        state = 128'h1237_fba5_a981_76c7_0100_3bf3_b92a_0d4d;

        #200;
        key = 128'h3dda_03e4_e176_3821_dbf0_1b14_5506_1a45;
        state = 128'h0dc6_167f_1f22_b194_cbc2_1ba5_6166_8dca;

        #200;
        key = 128'h7b23_eac1_8036_c91b_7dd1_dbb3_5fbe_cfac;
        state = 128'h405c_80df_ce18_e1ad_4be9_5a2f_5684_4e68;

        #200;
        key = 128'h6850_dcba_2706_1087_54e3_80dd_18fa_bc73;
        state = 128'h99fc_d1e1_5c7e_69a2_5810_12d8_1a43_54d5;

        #200;
        key = 128'h06d1_6dc5_16ed_3d69_e37e_2e57_f023_af4f;
        state = 128'h90f1_b02b_634a_8099_ecb9_ab8e_bbd5_1003;

        #200;
        key = 128'h0ff5_c8fb_439e_96b9_696c_9577_3cdd_b285;
        state = 128'h578d_7a80_6d6e_aa36_64c1_c927_d45b_cfc3;

        #200;
        key = 128'he14b_6e7d_2f53_9af8_5b01_68df_1342_df0c;
        state = 128'hd9c2_f493_21fc_d3ad_8881_1e3d_cc8c_dcb0;

        #200;
        key = 128'h3abf_b7d2_d38c_cb92_05f8_2ef7_49ff_7f03;
        state = 128'h53f7_4c1a_3552_6cbf_0f54_e27f_3d19_42dc;

        #200;
        key = 128'h58a9_12ac_e445_b341_f193_b8bc_2c33_7245;
        state = 128'h0386_0853_6ce9_3bcd_c1a6_2b34_02d8_5917;

        #200;
        key = 128'hdc9c_384b_fcdc_cfa4_a31f_87a6_838e_aca7;
        state = 128'h1cd3_7fa4_8f3d_4c23_746b_921f_74aa_7331;

        #200;
        key = 128'hf471_439b_159b_895d_60dc_aa8d_fff4_6742;
        state = 128'hc0d7_a5da_3dce_4ced_721f_5a22_5aca_28e8;

        #200;
        key = 128'h84f0_9b37_749b_2b86_c752_ca6e_2610_65fc;
        state = 128'hb0ec_19b9_a75a_40b5_ab7b_0e6e_252f_ab3c;

        #200;
        key = 128'h9637_76a9_9b08_11f9_8ebf_2977_a55f_4586;
        state = 128'h3fdf_6303_d1f9_6859_2498_756d_be19_1b77;

        #200;
        key = 128'h5e31_ef16_82b9_8c93_2355_705a_fa2c_32e0;
        state = 128'hf0b6_786e_27d7_61fb_9500_d773_0fa7_e0a7;

        #200;
        key = 128'h4ecc_d2b8_6dd0_096c_aebe_77c0_c4f8_d191;
        state = 128'hfed3_f299_7dcf_d158_8249_60e2_3fad_62cd;

        #200;
        key = 128'h4af4_3c21_08be_d799_4acf_66bc_1057_0a45;
        state = 128'ha16e_4aeb_09df_f981_0b88_861d_1616_a5e7;

        #200;
        key = 128'hde78_c8e4_1436_8b07_6ca3_a06e_04b1_4550;
        state = 128'hb1d4_e2e5_c4d1_8503_dc88_2fcb_a4fa_2e76;

        #200;
        key = 128'hc59c_fa6c_32ca_bc5e_ad62_a218_a5b0_7a0b;
        state = 128'haf4a_27e0_f7c8_b15a_e5e6_79df_201a_5132;

        #200;
        key = 128'h5f3b_f440_d436_480b_45a5_d277_27df_7961;
        state = 128'h82b2_e2ce_ff3e_4aa0_6a5e_c342_1f7e_8344;

        #200;
        key = 128'h40a6_9bb5_e503_05e2_1c51_c955_e34a_1aee;
        state = 128'h9b40_4227_c7d4_b346_9122_25c6_097c_db73;

        #200;
        key = 128'h5c1f_eb87_ce90_6abd_3199_a4d7_9bf2_a8a1;
        state = 128'h390e_3e66_7987_5046_f05e_c1c3_5fd4_4e68;

        #200;
        key = 128'h0097_b3b8_faa1_62f1_a4dc_8302_3e65_60b7;
        state = 128'h7f1d_f992_5ef1_463b_2b87_7614_553e_fc3e;

        #200;
        key = 128'hab88_bb40_56ee_cd8b_d565_4a82_e634_e9cf;
        state = 128'h19f0_f10e_2ecd_0b21_25e6_0bc9_b527_b635;

        #200;
        key = 128'h5f88_ff1a_af9f_1e06_6e5a_1e15_0065_fc66;
        state = 128'h9290_7aac_eabd_6307_c518_cead_d6f7_1fa3;

        #200;
        key = 128'h2e4a_20fb_8feb_8189_f14f_4d70_d2d3_45eb;
        state = 128'h276d_044b_be30_7d9d_0802_51d1_dcfa_eedc;

        #200;
        key = 128'h7975_6435_aac3_873e_1be3_dd27_a18b_592c;
        state = 128'h3dd2_cf16_e7f6_6ad5_654f_8ebc_bc84_0fc4;

        #200;
        key = 128'h95c9_2101_d4e3_b237_e4b7_4f5e_c32a_6358;
        state = 128'h3e8e_7b2e_2573_401a_085d_9722_16d9_67ff;

        #200;
        key = 128'h61bc_fbef_b7d1_ad6b_0ba5_4964_3798_ffc8;
        state = 128'hd9ad_862f_5894_ce79_7bda_fc1b_a55a_1503;

        #200;
        key = 128'h2248_21f1_6004_eaf9_d322_a384_83b5_9e2e;
        state = 128'ha88b_f14c_bd37_9adf_9017_db6e_2fad_e87c;

        #200;
        key = 128'hcb23_fc10_0ad8_1d17_6111_e603_47fe_b6e4;
        state = 128'h3a4e_2548_9502_6fe0_2ef3_2a21_0265_5852;

        #200;
        key = 128'h4d4c_40f9_b3e8_643c_b9a3_d69b_8ab3_1ba5;
        state = 128'h6565_02b1_a45d_e3c7_0f13_d09b_acaa_2600;

        #200;
        key = 128'h2543_b652_1997_b374_3604_49e5_9bfe_cbb5;
        state = 128'h2b68_8970_a852_2159_1461_46da_36cb_ad0b;

        #200;
        key = 128'h42ca_5b1d_69aa_c02f_783a_b682_34ae_5fab;
        state = 128'hfd5c_507d_6820_60de_1c09_1ea2_81ab_e3ea;

        #200;
        key = 128'he121_7e40_1862_961f_7913_ffdd_3edd_9ac6;
        state = 128'h5d17_f221_9384_ae08_1994_2dc8_ebc0_2502;

        #200;
        key = 128'hfa2b_6fc3_a9d7_b514_e247_7a0f_5f96_f59e;
        state = 128'h1570_56d1_a4f5_dd23_928e_a627_baac_af29;

        #200;
        key = 128'h9da2_af17_6caa_1b0b_1b46_617a_5ba9_9844;
        state = 128'h992b_012e_5428_30e7_55c4_078a_0ac6_065a;

        #200;
        key = 128'h9527_d04d_a0a9_18d9_6088_fa41_ce0f_850f;
        state = 128'h2024_8a21_613d_3ad5_734c_4757_4261_4b6e;

        #200;
        key = 128'h886d_7b3e_28b5_54de_a70f_ca91_9ef1_e061;
        state = 128'h01ad_c1c8_b1e1_0e13_ad67_eaa0_58a9_2910;

        #200;
        key = 128'he369_9f2f_67fb_ba02_7969_16f1_617d_0dd7;
        state = 128'ha23f_25d1_9f74_bb4b_cfa2_af54_2875_7d08;

        #200;
        key = 128'hcefa_44f8_0ad2_0c04_6a2d_98ca_e2ea_6400;
        state = 128'h7d46_bbf6_57c9_d159_04d3_b39c_4ffa_274b;

        #200;
        key = 128'h527d_f665_8f8a_0e48_4788_fba6_86cb_538e;
        state = 128'hf915_6e29_9499_1ee1_e519_2f1a_0fb3_b933;

        #200;
        key = 128'hab36_3739_dfcf_cb42_a203_5030_07f4_e8f2;
        state = 128'h0f82_6e62_859c_b708_137b_42ea_6367_bbee;

        #200;
        key = 128'hca8d_821d_9ef9_c5c6_da2c_7d18_1605_49ca;
        state = 128'hcd1f_7e0d_1547_96ca_d5f5_e43d_0365_2058;

        #200;
        key = 128'h384c_a6c2_ed5f_80c3_5ed2_05fd_83d1_5127;
        state = 128'hcd1b_e575_95b5_b1e2_06a3_9842_a91f_fa28;

        #200;
        key = 128'h7198_11f1_c561_9567_0747_2812_4cbb_abe6;
        state = 128'he595_4587_4f95_edb3_a83f_655b_663f_07d5;

        #200;
        key = 128'he0a4_2bb1_3470_500a_06d4_6faf_294c_eff7;
        state = 128'h947d_3b16_8294_dcbc_d11c_839f_5a20_56b7;

        #200;
        key = 128'hcc0a_08ba_bf3f_bfff_892d_32e8_5ded_9d9d;
        state = 128'h8da7_1735_c478_dced_d767_62ef_e347_c3d6;

        #200;
        key = 128'hf38e_0414_462c_af3f_b5a4_b26e_c3a2_7224;
        state = 128'haa71_e7dc_8d67_8e14_3ffa_a74f_bb02_9d5c;

        #200;
        key = 128'h280e_f6eb_48b1_5ca6_891b_4144_b2b7_71ee;
        state = 128'ha7f5_2cc7_a5b1_05be_aeee_4eac_fcff_f8a8;

        #200;
        key = 128'hef6a_ae0b_932a_3517_7e47_b9a3_bbfe_621c;
        state = 128'h3270_dc5c_ea2c_4fb7_381a_dc6b_23b8_5fe0;

        #200;
        key = 128'h0939_bd65_35ed_36bc_296a_4e15_5a97_f1da;
        state = 128'h9b20_2058_9779_ee27_632f_e3e1_ad2b_9c34;

        #200;
        key = 128'hba37_4f0e_b30b_e390_a790_10aa_e77c_70b1;
        state = 128'h7db9_6f52_c801_2abd_159e_b4dd_fb68_199d;

        #200;
        key = 128'he6e8_8b75_19a9_d3e3_f308_d83b_6f73_a5bf;
        state = 128'hce18_7323_4cac_4630_1685_5f09_5406_29de;

        #200;
        key = 128'hd4c3_c413_c5b5_3401_3815_23b8_7acd_36ed;
        state = 128'h7e6d_0606_8a9a_4b34_ed65_9ebc_6cf9_c370;

        #200;
        key = 128'h706d_c67e_0996_309c_9a49_8cf9_8052_26ee;
        state = 128'h679e_8d71_4bac_97dc_6f2f_2536_a3cb_84b5;

        #200;
        key = 128'h9f73_4ee7_9a3a_0f60_af59_3982_5017_8e4d;
        state = 128'he66f_5428_a2f9_5b71_64ce_72ff_6d5f_d89b;

        #200;
        key = 128'hd6db_2b56_7b82_7517_ddf0_962e_9877_0fbe;
        state = 128'he6f6_abc9_dadb_cfcd_bab6_f7a3_77f6_5387;

        #200;
        key = 128'h3cde_3bed_90b3_c68a_542c_cbf2_9fc4_31c0;
        state = 128'h1e00_fc5d_6a3b_a644_1609_2121_a76c_f262;

        #200;
        key = 128'haae8_4041_30c6_8309_905a_50db_422c_f4be;
        state = 128'h9504_1f39_7de5_af88_aa0b_b054_0c8b_3ebc;

        #200;
        key = 128'hf5cf_ceaf_834b_74bf_ad1b_9e95_aeab_9cd6;
        state = 128'hd532_9bbb_e5f3_b117_48a7_4ccd_c1ca_227c;

        #200;
        key = 128'h19a4_8b1f_4e8b_c3aa_9ff8_6fdb_d399_319e;
        state = 128'h4915_d859_f436_639b_07a8_5453_94ba_4039;

        #200;
        key = 128'h3ee9_d669_45bd_d36b_6d12_097e_3de1_4ee3;
        state = 128'hefae_afdb_bae4_601c_e720_115b_61b4_0a6a;

        #200;
        key = 128'h7134_4eb7_72c7_da7e_95a4_469d_91d4_8770;
        state = 128'hbd87_f25f_07c4_01f7_d573_1037_e438_47f8;

        #200;
        key = 128'h9870_1411_662a_f9f1_a02e_32ba_bdf2_f52c;
        state = 128'hb65b_495f_c71f_b168_ca2b_4ddf_56a8_feb2;

        #200;
        key = 128'he88e_63ce_3c57_8923_6617_0573_4c37_1392;
        state = 128'h08da_12fc_df1f_d04d_417c_9563_a976_8c9b;

        #200;
        key = 128'h97fc_63ea_d0f2_e928_66d4_3ccb_17a2_2e0e;
        state = 128'h237d_b939_9822_011f_80e3_3b34_8c57_42cb;

        #200;
        key = 128'h88a0_862f_da17_3cba_9b9b_d5f9_ddec_69c6;
        state = 128'h3d7b_b7c6_1870_20bb_4f67_1793_6e7f_11fd;

        #200;
        key = 128'h0bf0_38a9_dddc_fb3d_d66d_8537_6ee5_ee81;
        state = 128'h19e4_e5e3_7af1_cc35_85ba_75f9_16d2_8839;

        #200;
        key = 128'h2a9c_c35f_7560_50a5_4dd5_d30f_87c2_6403;
        state = 128'h28fd_2533_2c65_7403_cd50_9af8_deb1_e864;

        #200;
        key = 128'h9167_b2db_5488_1e44_5d86_7fea_fbc6_d8f6;
        state = 128'hbb05_1bed_edad_1b7a_07f8_7a82_8749_7a0a;

        #200;
        key = 128'ha727_c784_ad4b_4ad6_5f1e_6a7e_c021_4e37;
        state = 128'ha2f0_b7a0_e71d_d62c_f46e_0b0a_038a_52da;

        #200;
        key = 128'h40fe_7f95_27d0_fe9c_c43b_1869_1f8d_1717;
        state = 128'h8734_0c68_398e_9bc2_1e72_c7bc_cfa5_04a0;

        #200;
        key = 128'h1bcc_99b5_4d5e_0cf8_4b0f_0ec7_d929_181e;
        state = 128'h46b9_f088_e719_c742_68a3_1e2a_dab2_2bd6;

        #200;
        key = 128'had0f_1702_408b_732f_a16a_1053_16b5_2919;
        state = 128'h7cc5_6f3c_75ff_184c_695a_1093_5a2e_a2e5;

        #200;
        key = 128'hb601_698a_2fb0_b534_2e00_da5c_96b9_7e91;
        state = 128'h076e_bd81_7a5c_bda0_8109_0a2d_919a_322b;

        #200;
        key = 128'h0f8d_fd6b_d09d_2eab_c77a_a597_35a6_c2fc;
        state = 128'h2d62_891c_c461_c79a_8c73_8437_66c6_b4f6;

        #200;
        key = 128'hbdf5_6f4f_2b7e_ad36_79a0_2cdb_4229_d711;
        state = 128'h8337_ec69_e059_a490_e5de_f0ef_5fae_c601;

        #200;
        key = 128'ha078_3f33_2f43_0a58_a3ab_3a11_2bff_d970;
        state = 128'he420_caeb_2c92_180c_9dc4_d773_403c_fba7;

        #200;
        key = 128'h4ce3_60f0_9035_aed6_ed32_46d7_c0f5_b4d9;
        state = 128'h789e_345a_f4e1_6d19_f1dc_d8e5_69dc_ddbe;

        #200;
        key = 128'h2625_46bb_086c_c174_a56b_f608_afbc_d3af;
        state = 128'hcf09_99d4_f832_498f_5731_39c3_aade_91f3;

        #200;
        key = 128'h68ac_a2bd_32d8_e8b5_bebc_a1a0_e024_6a20;
        state = 128'h60e2_971a_08f7_3b0e_cd5b_313c_fdcf_58bb;

        #200;
        key = 128'h9ed7_e125_fc5d_a9a5_c3d4_2e6d_dd2f_20c6;
        state = 128'h376c_a172_b3e5_4d39_4f6e_6621_c553_da64;

        #200;
        key = 128'h21b8_3056_4702_6ae8_e509_fa7d_4f09_40ce;
        state = 128'h6576_2958_4031_7d9a_cf4c_bf62_f2a5_ebc8;

        #200;
        key = 128'hb5bf_6944_836c_0ffb_a704_e0ce_3a0c_b5e1;
        state = 128'h8cad_67ce_df42_a732_b6c2_9bd4_0494_7d34;

        #200;
        key = 128'hc58a_457f_6a40_ecef_14a2_9629_5bde_3e97;
        state = 128'h4dbe_01fd_26da_4461_2957_c91e_e9d8_89f5;

        #200;
        key = 128'hb246_ae0c_1f4c_1137_aaf7_a789_476e_c888;
        state = 128'h9761_15e3_f356_2d36_3d47_a2e3_cc79_2967;

        #200;
        key = 128'hbe48_addc_3dcc_bf59_574f_b2b7_cc9f_d1b6;
        state = 128'ha111_6bc2_9eb7_112c_bfb9_77ae_412f_1ad2;

        #200;
        key = 128'h0982_01d4_15dd_5613_0e12_1e4d_831c_cc57;
        state = 128'hfd80_277e_f8c8_0e29_24b6_c98e_1bf6_988e;

        #200;
        key = 128'h3d84_af8f_30ed_3432_62b6_f36d_c26f_1b92;
        state = 128'hfcd8_e507_52a8_7598_a910_6464_4b25_b76d;

        #200;
        key = 128'h1e94_90df_8627_9b08_68de_4ddd_27a0_770b;
        state = 128'ha656_9cf6_a853_496c_fe6c_6604_3032_1b13;

        #200;
        key = 128'h8734_8184_5064_6dda_488f_cc92_08f6_7286;
        state = 128'he282_0dea_a091_74a4_0771_bea7_020d_249b;

        #200;
        key = 128'h68be_c2d4_1ee5_8da7_21bb_5fba_6a04_d147;
        state = 128'h7320_345f_e988_cb94_121a_949f_c5c4_9881;

        #200;
        key = 128'h1ed4_c280_0435_73ef_954b_cfa2_4c28_babb;
        state = 128'h334e_9c97_5175_aafa_1fdc_f171_5928_9234;

        #200;
        key = 128'h334d_b6c5_ff6d_8e74_86d0_b7d0_304a_e457;
        state = 128'h9c0c_ff07_620d_6fbb_af8f_c11b_d4e6_a9ad;

        #200;
        key = 128'h6806_4676_90df_e53d_1552_09db_36cf_0c74;
        state = 128'h177b_e883_2bfe_4398_c3e5_3dc8_a88e_06c5;

        #200;
        key = 128'h2195_604a_eac8_1a07_1a37_4dd3_b4e6_7813;
        state = 128'hd2f6_793c_f430_b245_c673_733f_078e_9bce;

        #200;
        key = 128'h0cb6_9771_ac71_5245_ff2b_d9c8_baf9_e522;
        state = 128'hd0c5_79be_4976_0025_02fa_5848_ce23_4b0e;

        #200;
        key = 128'h6d41_eb47_bcdc_9b26_6b15_1101_2af4_1ca6;
        state = 128'h97b5_157d_4549_4292_f158_6783_cfae_07b3;

        #200;
        key = 128'hba10_ec67_3c9f_d2bc_1018_b958_8776_2e5d;
        state = 128'h582b_5c6c_a913_7641_ebaa_94b1_2228_b7de;

        #200;
        key = 128'hb5c9_0550_2677_12af_205e_6b0f_5673_788d;
        state = 128'h0e98_2545_78a1_447c_5fd1_9342_1f75_623c;

        #200;
        key = 128'h266c_80d1_43bf_cc21_f92e_716e_ba1a_f9eb;
        state = 128'h60af_ae8d_d918_9170_d990_9105_5d94_eee6;

        #200;
        key = 128'hcef2_684d_abbd_99c6_f9ee_8dc3_4969_bb60;
        state = 128'h9b99_8a05_1ec3_9516_f2ef_c713_f81b_207f;

        #200;
        key = 128'h8baa_ecaf_274c_fbdf_eee1_e73e_bdd0_1303;
        state = 128'h8b4f_73d9_601e_aa6d_272b_1b60_2918_e2ab;

        #200;
        key = 128'h11f0_affb_6f6c_f384_c73b_8c9b_e7af_8656;
        state = 128'h5e39_2e69_77fd_6f47_2d19_dfe8_ef82_77a0;

        #200;
        key = 128'h8b9d_b7de_e95f_0743_ea0e_9807_0e6e_3187;
        state = 128'h5a7b_246e_946d_1374_ccd4_c41b_7264_463b;

        #200;
        key = 128'h50c4_35ec_960e_d3e7_b728_ab0f_6969_1f1f;
        state = 128'hfdbd_8e25_4975_2525_7824_c00f_2d8e_5eb3;

        #200;
        key = 128'hb707_4ba6_a7ab_fb79_3065_a186_30a6_2552;
        state = 128'he296_782b_db96_8778_cad4_dc68_8a35_221e;

        #200;
        key = 128'h6971_779e_f680_b330_578d_c54c_a31d_3193;
        state = 128'h6956_16f4_9693_41a9_5c7c_b79d_0c8e_6592;

        #200;
        key = 128'hdb7e_7348_3f84_36f5_d9af_a1a0_ea32_5140;
        state = 128'hbdf1_4ccb_d071_4885_8675_764a_e246_7581;

        #200;
        key = 128'h1ed9_c7f3_b9c7_97d5_8675_40ef_0561_d46a;
        state = 128'h4569_4a47_c43c_a943_9303_01ec_339b_4545;

        #200;
        key = 128'h43ca_2865_ffe4_823a_8481_0526_c7a7_98ab;
        state = 128'h0268_4d13_fece_24ee_0b2e_5cc7_ef25_f1eb;

        #200;
        key = 128'hfaff_29d4_9d08_cb10_0f91_8128_624c_3bd3;
        state = 128'hd184_4039_46f9_cd43_69b5_0ee3_bfe9_a30c;

        #200;
        key = 128'h618b_770f_0098_4ba7_bf83_e42b_3307_5a0f;
        state = 128'he69f_c59a_8bc8_af15_a3e1_ec7b_3e2b_8bc0;

        #200;
        key = 128'hcf2c_887f_da6a_b03e_6833_dc71_f65f_2918;
        state = 128'hb6a7_7025_2cad_8904_4709_6bdd_3347_e933;

        #200;
        key = 128'hf4c8_58f2_cd8c_5367_aadf_7954_6700_0f11;
        state = 128'hf180_ae65_11bd_7960_2d3c_0a5f_207d_ce10;

        #200;
        key = 128'hf825_719b_92e7_8a92_97db_4531_0758_e024;
        state = 128'ha1cc_aeaf_f133_c5cf_3cc7_3e55_3844_1d74;

        #200;
        key = 128'h4175_11d0_1c66_06b3_17f2_e245_837a_1837;
        state = 128'h75bd_e33d_c5d0_5df7_79c3_52b4_0932_7d11;

        #200;
        key = 128'h8a18_f377_ce19_4b58_8561_4ee2_5ec7_cda9;
        state = 128'hef32_5789_edbd_dda1_3f5f_4f2f_8773_c9fe;

        #200;
        key = 128'he6a6_fe2b_7196_56a4_5860_82b0_c646_a9ba;
        state = 128'hf6b1_de12_a2de_b97b_13d7_83cb_f1b5_e931;

        #200;
        key = 128'h0c9c_0b1b_5d3b_8be2_5604_534e_0271_7ab3;
        state = 128'h4fe9_7a5d_c459_aa44_83f0_97c8_4737_c206;

        #200;
        key = 128'h22d6_f22c_6be3_5e84_1bd1_ec6f_de1a_bc3f;
        state = 128'h8cb8_183c_6121_1824_4e6f_d95f_b73d_2851;

        #200;
        key = 128'h9614_8ee9_f283_8f26_2f7a_bbb2_d187_bb42;
        state = 128'h2489_0ab1_d6e7_a9d2_bd5c_60dd_acd5_1d5e;

        #200;
        key = 128'ha55f_d3c8_b980_f450_34e5_c07a_b939_f2a9;
        state = 128'he70b_3777_ff01_131c_2d1d_16e9_1723_c8c6;

        #200;
        key = 128'ha794_7b7a_cf26_b618_09b7_b22a_97bd_ed18;
        state = 128'hd2af_d6b8_e761_3c58_4722_628f_cee1_155d;

        #200;
        key = 128'hedbc_ecf1_6456_4d69_dfac_705c_5b26_80b3;
        state = 128'h6038_2adf_f13e_5e32_ce3c_e2a4_38f6_a8d6;

        #200;
        key = 128'hbb5e_1060_b0bf_dda5_d2a2_8527_714f_18b0;
        state = 128'h455a_6c22_4e9b_4098_2734_cf9c_7163_6bb6;

        #200;
        key = 128'h1880_dd1e_c03f_018a_448c_cff0_a4b5_53c4;
        state = 128'h7c23_484a_8341_66a2_5317_aa9a_d91c_5bd2;

        #200;
        key = 128'heec8_945f_c90d_b072_abba_3926_5438_712c;
        state = 128'h79d1_a5ec_6459_a000_db0e_d350_56be_4bda;

        #200;
        key = 128'ha43b_2159_6740_693c_7462_1a6d_3bc3_e93e;
        state = 128'hb7ac_447d_494b_e113_906c_a15d_1aa0_090a;

        #200;
        key = 128'h9a0f_7aaf_72cb_249f_f28e_3a61_eb0c_f523;
        state = 128'hb1ec_48ac_3d5e_e3f0_545e_f5a8_8a1f_e47a;

        #200;
        key = 128'h4c08_8c2d_919b_1b24_5243_f21c_cede_dff2;
        state = 128'h5827_8f06_b3d8_24e4_836b_ef1d_6431_a2d6;

        #200;
        key = 128'h2e5a_7353_4105_a7b8_a2a9_0319_5122_755c;
        state = 128'hec38_9d0c_7034_50d2_3bfa_8494_e262_6686;

        #200;
        key = 128'h399e_b7b5_2828_9136_3b2a_b188_281e_53c5;
        state = 128'hf7e2_0136_c36f_8658_0f59_40d8_c748_88b4;

        #200;
        key = 128'h3943_c5c3_a26c_a4fc_3bcb_3e43_ea68_d320;
        state = 128'h923b_beaf_d4be_40a0_5116_4958_1456_b930;

        #200;
        key = 128'hc4b7_009b_49f4_8cd2_b2b4_63bb_1a62_1c45;
        state = 128'h2d83_38a5_87fa_c2a8_abaf_527d_f5f5_fca7;

        #200;
        key = 128'h393f_a32b_c5d5_788f_2094_c663_48f9_a492;
        state = 128'h56a9_c14a_4bde_40e3_369e_0990_83c7_3d9b;

        #200;
        key = 128'h819e_2dd6_f4d9_2358_8c94_4693_6951_3955;
        state = 128'h5c0d_91d7_67e0_af31_c4fb_d234_8133_3090;

        #200;
        key = 128'h8055_a906_7259_3b0c_c7b5_960c_9480_13f9;
        state = 128'h306b_22c6_76a9_1182_de13_6da2_9a47_c69a;

        #200;
        key = 128'h4f5c_7467_fa9f_3e42_d663_fbdc_a18b_1757;
        state = 128'h34ae_9151_6f58_a011_3de6_d921_27f9_326f;

        #200;
        key = 128'hd76e_bacd_975b_d714_11b9_b991_bcd6_b346;
        state = 128'hf117_1d38_e25d_cc54_302e_156b_f508_6a5d;

        #200;
        key = 128'h51f3_467d_6d3b_df3a_8b6c_3c4d_997b_6ae9;
        state = 128'h8f3f_f06b_a18a_9018_285a_f4be_f376_f204;

        #200;
        key = 128'h6a51_6d76_5597_dc06_00a0_1301_4852_e5ab;
        state = 128'h50ed_ea99_9d4f_f09f_dde5_3c87_727a_1e0e;

        #200;
        key = 128'h5af2_b2cf_5122_0f40_12a7_df3b_7fa9_8c28;
        state = 128'h4396_dcf3_bd74_6c24_e5ee_1d24_db81_8b7f;

        #200;
        key = 128'hc765_1ef1_061a_ebe5_dfdf_7c78_7960_3777;
        state = 128'h7842_e979_6586_97ff_4312_5342_bf90_c486;

        #200;
        key = 128'h145d_5138_6d01_e6c0_61f3_456b_70b1_f3cd;
        state = 128'h9bd0_bb0d_b2ba_eff1_9142_104a_6168_8ff0;

        #200;
        key = 128'hbe7e_b268_290d_6d5d_549d_9bdf_f96f_a71d;
        state = 128'h7539_fcde_4834_9834_f34a_3176_ef73_16ac;

        #200;
        key = 128'h610a_15ab_ee23_3274_e688_db0d_dceb_62d8;
        state = 128'hda2e_afa8_30f0_d7fe_964c_32e4_cea3_1e76;

        #200;
        key = 128'h41bd_7e99_6e5c_f201_24a3_374e_c9e6_02d9;
        state = 128'h1e65_d9a6_7a33_26d2_bee3_52ff_51f1_e33e;

        #200;
        key = 128'h5603_d964_473a_0f84_80ff_0f9c_a66f_688d;
        state = 128'h4cef_ea24_b405_9ba1_9ac1_42fe_6229_81b2;

        #200;
        key = 128'h1332_59be_0b76_eeab_c885_92f7_7a29_3d9d;
        state = 128'hda54_4af6_bbce_9db8_7c52_8498_47f8_ca4a;

        #200;
        key = 128'h76f0_bcc3_1ec8_0be2_8eba_2c7d_ba0f_e867;
        state = 128'h9740_e3ec_20e0_6502_9b9e_9d70_7f40_b445;

        #200;
        key = 128'h0488_5b48_2452_1cea_9e53_9417_6938_3334;
        state = 128'h92c3_28ff_ef5f_75f4_3c85_200a_888c_cf24;

        #200;
        key = 128'hb507_20a5_3918_b8fd_5b2a_cccd_967e_c7e2;
        state = 128'hf2ec_2d1b_029d_9dc7_4257_2869_9ed1_6cf0;

        #200;
        key = 128'haa4d_aeb7_2181_0d97_1f47_94e5_4ce0_41e9;
        state = 128'h2d25_6f1c_0d12_e2b8_4f3f_3561_7eb3_33c4;

        #200;
        key = 128'h5915_f6ad_dc33_2025_d4f3_f56d_2ec0_fc2b;
        state = 128'h0394_5118_471b_b0fb_df39_8bf7_1878_f9e6;

        #200;
        key = 128'hde72_e84f_1500_a571_8e73_6e0a_e914_690d;
        state = 128'h7619_e651_f03e_7ab6_6c0d_d05b_1e90_4721;

        #200;
        key = 128'h97f9_ce20_90d4_438b_cd78_e4be_caf8_a89c;
        state = 128'h227f_1dcb_349d_2eac_eb71_a10e_d5e4_4c02;

        #200;
        key = 128'h810c_3cf6_26f8_07a7_ea7d_0b27_c985_e001;
        state = 128'h0184_6ec0_2706_1509_4c3b_eec6_6fcc_fe62;

        #200;
        key = 128'h2d00_6b47_cbb0_832c_9189_bc8c_e48f_a110;
        state = 128'h1b9f_e020_5649_a174_db96_8c5a_c29c_aec6;

        #200;
        key = 128'h749b_0b7a_04c8_28a3_9bea_52a0_3985_042b;
        state = 128'hf39e_0537_18da_5ac1_29ec_90da_c923_e3e0;

        #200;
        key = 128'h22c2_eb79_9e9e_9572_acdc_edd0_1872_a2af;
        state = 128'h157b_781d_1c85_f322_eae3_c8ff_9008_00a2;

        #200;
        key = 128'hce88_72d8_79e3_8cc0_c8a4_8645_023b_fc85;
        state = 128'he5f7_e48a_944b_9c9d_1b70_0e99_1b65_75aa;

        #200;
        key = 128'h83ae_a402_c59a_3378_6241_6ede_716a_feba;
        state = 128'h4ed3_727e_bc67_19d3_1f82_41e8_3507_9166;

        #200;
        key = 128'haaf9_db18_eaec_eebb_0bff_d40d_88d0_500e;
        state = 128'h5b0c_7c38_de44_b8b0_e1b2_a77e_e606_696c;

        #200;
        key = 128'h82fd_66cc_4df2_a069_862e_c535_847e_1336;
        state = 128'hff8b_cefe_a266_a6fe_3aa0_2bf2_2c70_2d6d;

        #200;
        key = 128'hfc90_78d9_0c0e_f5c1_0d1f_3064_f3b9_1a9a;
        state = 128'hb94f_ab76_cf09_9ad5_d7fb_e545_2aea_4e3b;

        #200;
        key = 128'h8087_e002_7ad3_6b55_3bba_dc94_7989_5f7a;
        state = 128'h3781_d762_f82f_6a42_0e94_2799_0f96_52a3;

        #200;
        key = 128'h5dbd_b773_8058_423b_141e_2b06_89fa_23f8;
        state = 128'hd4e1_7562_175c_5dd2_c82e_b6ea_cfc2_e3cb;

        #200;
        key = 128'h74ee_4713_179b_2e47_b776_3bfa_0672_8bad;
        state = 128'h432e_c8ca_ff08_53e2_28bd_3ee2_0d68_ffb8;

        #200;
        key = 128'h9200_c965_a239_cf9a_8a78_9896_eed7_6c76;
        state = 128'h79ea_2d1e_1eb6_0dac_8c6e_f054_c968_05f0;

        #200;
        key = 128'h315c_955d_c53f_98f5_7452_1e6e_82ba_f1a9;
        state = 128'hc7c2_60a1_03df_c0a4_a228_0a48_5148_89e5;

        #200;
        key = 128'hdd3b_88e4_6982_8731_76c9_570d_2366_4513;
        state = 128'h1175_0830_1742_21f7_cfbf_9441_9e94_03ce;

        #200;
        key = 128'hdb17_a312_51ac_3e17_1e38_473e_e2cd_2491;
        state = 128'h87c3_6741_c9fe_983b_cc7d_2d77_15ef_ffd1;

        #200;
        key = 128'h17d4_7b04_dff0_76ce_70ca_1ab9_fc8b_657a;
        state = 128'h50ce_6d72_af21_a0eb_32ed_b606_28a4_1f79;

        #200;
        key = 128'h9018_6acd_1a45_3a94_6347_69fc_e225_beaa;
        state = 128'hd9b5_8b16_7cfe_5b09_42ec_fe81_5d21_53cf;

        #200;
        key = 128'h81e5_08c2_65d8_0f52_be7a_ced9_7d6c_a432;
        state = 128'h3686_a745_4e58_6a55_146c_7521_8ce9_a857;

        #200;
        key = 128'h4aaf_8e64_1258_f8c0_900e_48da_56f8_d727;
        state = 128'haa7a_d94d_7e22_618b_7215_82d1_627f_7e71;

        #200;
        key = 128'hb663_8512_b2d0_9e05_8a0a_be06_83aa_3c34;
        state = 128'h00eb_4c8d_6555_fcda_4ac0_e354_f054_0660;

        #200;
        key = 128'h64c2_283a_da0a_5ebb_a4a4_92da_6e3e_2e66;
        state = 128'h59ce_0908_17af_f510_d057_523a_b191_1fb4;

        #200;
        key = 128'hf367_a08a_720e_7069_45d3_8adc_c568_cf29;
        state = 128'hb764_bd04_398b_5b45_401d_662b_8126_5cd9;

        #200;
        key = 128'h1832_0e1c_922b_6bad_eafa_724a_d91e_1174;
        state = 128'hd3a1_7300_3f1c_cca1_4114_736c_5608_65e6;

        #200;
        key = 128'h39ca_842e_ce3e_611a_f01d_e477_ea6f_289b;
        state = 128'h2e1c_fff3_9acc_ce8c_bc57_2c6e_a8b4_72e8;

        #200;
        key = 128'h43d1_2508_308a_c8f1_f1c5_2690_2d64_0bc6;
        state = 128'h1fb4_4fcc_7efb_9572_ce5f_4034_2c0e_ad30;

        #200;
        key = 128'h1c31_0e9d_011d_6dde_56f7_2813_110f_2c8f;
        state = 128'hb740_71e9_f8cc_aca5_731a_b9a4_3113_5ae3;

        #200;
        key = 128'h8ba5_3d11_c0f7_9247_6f21_5504_c9be_5069;
        state = 128'h3d73_9c1c_3e5f_f846_288e_2f84_5547_ed52;

        #200;
        key = 128'h8ce3_bea8_3f76_f2ae_0c72_43c2_d923_c9a9;
        state = 128'hb99a_e0f0_71c8_cab0_3bea_b8cf_62e9_d50b;

        #200;
        key = 128'h9e57_fdc4_f7d5_a2b1_05d0_fbc1_db77_c891;
        state = 128'h8f27_b641_53fa_a60f_04e7_79e3_1331_cb98;

        #200;
        key = 128'h1071_310b_f3e7_e801_c94d_3f51_e88b_47ea;
        state = 128'h2d14_c336_7475_511f_bc97_751c_58c8_bd1f;

        #200;
        key = 128'h1bcb_361d_c54c_7dc3_cf38_c602_e2be_2bb7;
        state = 128'h71bd_7004_1391_332b_f945_5528_a8e0_3417;

        #200;
        key = 128'h37cc_1c76_2a65_9b25_bc74_5fc7_71eb_047a;
        state = 128'hfd30_04f5_4dc6_ed01_fd5d_7fde_6f36_0a7e;

        #200;
        key = 128'hd23c_54c5_2a37_6df2_1c0e_0d35_c661_7833;
        state = 128'habe4_8ca6_0d58_ff6d_d858_cf51_3d51_a597;

        #200;
        key = 128'h6ad3_5ea8_94f1_4859_2048_8178_fca6_4255;
        state = 128'ha76d_deeb_0c84_2ae5_1a0d_a779_b329_ff35;

        #200;
        key = 128'h607f_be93_c604_c677_9ffc_8b7a_0201_d8ed;
        state = 128'h6e68_8731_6eed_be5e_abcc_6d1c_4b49_3030;

        #200;
        key = 128'h9cb2_a884_8a8d_31cc_254d_e96f_14e5_a27c;
        state = 128'h3d38_f2d6_5136_0270_3a36_1b2b_1ab9_539c;

        #200;
        key = 128'he6b8_634a_da8f_f114_0cf0_206b_f869_33c3;
        state = 128'hf5c2_1791_6bd3_a9ba_b4ee_b890_18d3_2221;

        #200;
        key = 128'h695d_b0bf_71ab_6c13_c908_68ab_f9dd_7993;
        state = 128'h2d0a_0c9b_86d3_7cfa_3d0e_1276_951f_65d4;

        #200;
        key = 128'hd6c7_a0af_72e7_2644_8437_0ddc_3138_8027;
        state = 128'hf9f9_326b_bf75_8baa_14de_6f5d_c8db_5028;

        #200;
        key = 128'h39f8_a404_1608_17c1_e59d_52ce_e9de_1582;
        state = 128'h80c0_253d_ae12_5d40_741c_89fd_2c74_d6ba;

        #200;
        key = 128'h02cc_f028_052c_f16e_5b17_0bca_6340_2a82;
        state = 128'hf41b_2d99_c61a_28d7_9f6c_0e63_7263_90a5;

        #200;
        key = 128'hbc03_80e6_4eea_01ea_7a5e_b9d8_177f_5f7b;
        state = 128'hf0cd_be21_a903_af25_5ee1_c961_d1e8_1ed5;

        #200;
        key = 128'h59e2_5192_acc3_e004_1436_436e_9bd3_164a;
        state = 128'h05a5_72dc_d677_42fc_05e8_d661_e68e_33c5;

        #200;
        key = 128'hfec1_c522_9de6_6ed8_9d86_de54_564e_738b;
        state = 128'h9ea6_cd3c_e3eb_d816_b176_54ae_e96a_e02b;

        #200;
        key = 128'h3750_e50c_1940_e25d_9960_4049_e1bc_1c5e;
        state = 128'h363f_c208_c9f4_75bb_f67f_cd8d_99b8_c228;

        #200;
        key = 128'hdb38_8f7c_1a3c_c0e2_8e56_64c0_51fe_4b1a;
        state = 128'hdb8f_b9e5_e6e3_c57c_7fd6_02ed_19b3_3219;

        #200;
        key = 128'h792e_bd9a_788a_5540_ca6d_ee2c_381b_70db;
        state = 128'h572a_f9c2_6ead_febe_b9ed_e30d_3c0c_43eb;

        #200;
        key = 128'h2531_4650_78c8_d62f_ddda_f25f_c2fa_135b;
        state = 128'h8f82_0c01_ae10_91df_c3a3_276a_56db_fc37;

        #200;
        key = 128'h624d_49f0_c003_98b6_dd57_359d_a63c_b873;
        state = 128'h52f0_ea15_20f1_d535_7712_ddf9_41fb_d7bb;

        #200;
        key = 128'h8f1b_7409_f070_d1b3_8a0a_6c16_9c28_a138;
        state = 128'h7919_f101_ba70_15b0_7b73_cad8_67f7_d95e;

        #200;
        key = 128'h6c88_b9f5_4307_45cb_398b_d54c_8f7a_18d8;
        state = 128'h485a_5d71_f6fc_d8db_971a_2d7e_aedf_182a;

        #200;
        key = 128'hcf6c_d384_4c4d_0d42_7975_e3f4_229e_f02b;
        state = 128'h94f7_1570_ed8c_5b46_89a4_ca58_0179_f771;

        #200;
        key = 128'h1e4b_5ca5_37f0_fdda_490f_f36f_d264_319b;
        state = 128'h1f73_8182_cb00_7214_999c_af11_7748_08c8;

        #200;
        key = 128'hab40_403f_98df_7028_88e6_9365_2606_fbc9;
        state = 128'ha5e4_97db_57b9_27fa_9efa_75b0_e8bf_4abb;

        #200;
        key = 128'hfad9_c49b_e357_f369_a614_cacb_4d03_8a33;
        state = 128'hd2d3_5ee3_593b_a526_e214_11e5_4ea5_5364;

        #200;
        key = 128'hb71d_9594_7397_36b7_03cb_57da_522e_c249;
        state = 128'hfdae_76cc_0664_ef4a_e1f5_4721_2f13_c320;

        #200;
        key = 128'h0828_c02c_9d7d_765b_6cca_1666_70ae_ef95;
        state = 128'h9893_b176_9241_e7bc_9aff_e809_b58e_88b1;

        #200;
        key = 128'h98fe_a449_dd9b_9f88_414b_41b0_5544_144b;
        state = 128'h197c_db49_ba97_21ad_5ce4_0704_2e5e_c3a0;

        #200;
        key = 128'h8958_5f92_1a56_3af5_22a8_f91b_b06c_b9f0;
        state = 128'hc247_3220_ceaa_f6ce_72a0_4923_4e62_ea6b;

        #200;
        key = 128'h66d9_8d94_5c32_0521_2731_81a3_6f28_5bef;
        state = 128'h8733_50ae_99ca_0697_646a_ff14_046c_9c76;

        #200;
        key = 128'h8b5b_3c10_eae0_329f_d2cf_d7ec_5b41_8077;
        state = 128'hebac_ab25_1668_dc16_21f2_ec40_8f6e_8eed;

        #200;
        key = 128'ha11a_fed9_1385_e824_5081_15f1_5cf8_24da;
        state = 128'h37ea_8bab_414a_15ce_9767_a929_0a21_268e;

        #200;
        key = 128'hf133_e6ce_6e7a_8236_bcc2_2d68_8497_3e04;
        state = 128'h2f40_59f5_c55b_3c1b_3def_0e21_df0e_303a;

        #200;
        key = 128'h1955_6429_e7d4_828b_abcb_c035_ff98_6407;
        state = 128'h7eb7_7636_78b6_6b3c_68a6_3f4b_ca1c_884d;

        #200;
        key = 128'h6943_404d_e871_2fa8_7a69_a2c0_f32b_e6cb;
        state = 128'h7db5_d705_8100_e9ed_7d3f_d95a_8973_50c6;

        #200;
        key = 128'he179_2e12_ae12_3380_4a84_9275_6689_7b55;
        state = 128'h7dc3_d710_4dd6_5e0e_8a4e_60e1_c0ca_82eb;

        #200;
        key = 128'h0adf_2a16_5c5f_ecdf_93ea_b0b4_6fdf_07e9;
        state = 128'hb04d_2bc5_aa9c_1b5c_bee7_0f0a_9e3d_e044;

        #200;
        key = 128'h5d34_f00e_6712_2312_ea17_af8c_d4c0_72ab;
        state = 128'hc00f_03bb_84b3_343c_2bfc_1552_4254_5a4d;

        #200;
        key = 128'h8cdc_df43_19aa_5109_4ba1_d8dc_095e_5588;
        state = 128'hb6a4_ba98_d463_c7b0_270d_a90f_6160_f3f5;

        #200;
        key = 128'heff9_a65a_28a0_741f_df50_4e94_10be_396e;
        state = 128'h37c8_f33a_7b05_172d_0328_ee24_7528_3035;

        #200;
        key = 128'h53c8_dc36_9715_acb7_f276_323d_96ab_a5b2;
        state = 128'ha2f3_2da4_86de_3f1b_e160_6552_d24d_5c75;

        #200;
        key = 128'h240c_ecae_29bb_a69f_e78a_edf1_8bd0_e902;
        state = 128'h58ae_1ea1_e690_cc7f_5635_5501_f691_dbc2;

        #200;
        key = 128'h74d6_8588_4055_d02a_f2bc_1140_e4db_87d7;
        state = 128'h6415_2dc2_30f0_0420_2359_6dcc_42df_1ea0;

        #200;
        key = 128'h898a_4641_543b_3f22_7fd6_48f8_c9f7_aa06;
        state = 128'h9aa0_4c78_0088_8135_9d01_cec7_5f36_afb5;

        #200;
        key = 128'h61bf_b468_4147_6a5e_7741_2340_a45e_42c6;
        state = 128'h29cb_e496_f162_e787_aa3d_022b_a624_40f7;

        #200;
        key = 128'h9e14_268f_9e2c_0950_fa68_ac63_3054_f8ff;
        state = 128'hf1e7_0bae_ff42_35a4_1e54_c8f7_325a_8a10;

        #200;
        key = 128'h26e6_c909_213f_70f8_7367_32ea_3e84_aecd;
        state = 128'h687f_6d7d_77e1_46a7_2f27_be88_6fb6_31a0;

        #200;
        key = 128'ha1bd_61f9_b1df_ad90_e492_dcfd_0848_73fb;
        state = 128'hbcad_1efc_2617_d79c_95e7_3956_2e66_9b52;

        #200;
        key = 128'haab0_992c_cce8_ec47_e4b8_0059_f748_8166;
        state = 128'h7d84_d3b7_0081_121f_d9f0_dc2f_ea4f_d18b;

        #200;
        key = 128'h5739_cfca_6da8_8626_dd33_1869_2706_85e2;
        state = 128'hb2c5_c6c2_f990_94c9_ea3a_95e2_077e_59ba;

        #200;
        key = 128'h711a_2d01_1145_619a_c7d8_045c_cd58_8447;
        state = 128'h9616_28fa_6a81_01c1_1903_d5c1_2108_3867;

        #200;
        key = 128'hf8e7_c901_c1fe_0f0a_21b4_e529_51b5_6f0e;
        state = 128'h964d_9b5d_b1b2_4fe1_6408_0a10_e500_75fd;

        #200;
        key = 128'h9462_6177_9ae8_f151_2cc5_bccb_df66_8973;
        state = 128'hae77_b469_badc_9876_a3fd_3252_72ef_faa7;

        #200;
        key = 128'h1df2_cfd2_946c_dfc7_77df_af5a_36bc_145c;
        state = 128'h49c3_5713_4324_e782_1071_2575_d7f0_5cbd;

        #200;
        key = 128'h678f_b779_6dc6_606a_6079_96f6_2db0_b2e2;
        state = 128'h4d6b_7b57_875b_9603_62cc_2ec1_494a_8f4c;

        #200;
        key = 128'h6182_6831_bea0_8d3f_3909_f16c_ad3e_441d;
        state = 128'hfaad_9cd3_5ebc_c2d7_226e_09ed_4844_bcf6;

        #200;
        key = 128'h94ff_f6fa_b46a_4526_6c56_37d4_03ed_55ab;
        state = 128'hc8ff_27b1_823e_c82a_5392_6b97_a5f8_7f5c;

        #200;
        key = 128'hec99_4dae_e37e_cd61_8917_b7f6_59ea_f7de;
        state = 128'hbf74_17fb_0e75_37be_b85c_6094_8d87_86f0;

        #200;
        key = 128'hf04a_59ec_27e1_edcb_2d89_1bee_a79f_6331;
        state = 128'h9557_61c5_6aea_4b5e_899b_637e_a147_6acc;

        #200;
        key = 128'h70a2_4cbf_3950_cc11_f705_e3e0_52a2_62d4;
        state = 128'hf7d0_1dfd_0a37_173c_4a00_3af0_7b00_e1a3;

        #200;
        key = 128'h05db_16d5_b570_a6a2_77bb_5d8e_b0f9_e7ee;
        state = 128'h2e27_62f9_93cd_7ffa_03f2_bcce_d574_570a;

        #200;
        key = 128'ha3f2_f2e9_6163_f7ba_7478_cc24_8687_3fb3;
        state = 128'h96c9_ebc5_80f7_45b0_f5e3_c0e9_9c4c_c5d9;

        #200;
        key = 128'hd493_215f_5859_b585_5427_de7c_46af_680f;
        state = 128'ha002_b0d9_c246_d6d4_9fc6_9d16_a3d2_632f;

        #200;
        key = 128'h4cef_afcd_33bd_9f3e_dad2_f943_a29c_3bf4;
        state = 128'hc1b0_0ab5_ad3c_2a2e_3546_5705_5453_db86;

        #200;
        key = 128'h941c_3d05_3fbe_1c72_ae13_6511_2bcf_074c;
        state = 128'h4e55_adc1_cd1a_d730_4da9_323f_e2ec_3081;

        #200;
        key = 128'hb7f7_347c_1595_1255_9e7a_c96a_2e7c_9e1d;
        state = 128'h6e1c_4db2_6e36_78be_0626_a5fd_17b7_de2c;

        #200;
        key = 128'h9131_1f19_e311_4792_eb31_6bac_48ac_0d14;
        state = 128'h9b00_ebd4_9ca3_54ec_fbbb_fa39_03b7_6ad9;

        #200;
        key = 128'hb05b_304f_039f_755e_9acc_c488_e171_c647;
        state = 128'h08c0_e2b8_1544_fec1_3350_5893_dd4d_fb45;

        #200;
        key = 128'h3d22_cf2f_615e_65e5_8a1f_3750_5603_8d6c;
        state = 128'hd81f_4df6_7c48_774a_fb0d_faca_d7ca_30c7;

        #200;
        key = 128'h87a3_4973_af51_8d27_f251_0fa3_3769_3f4a;
        state = 128'h66c1_e915_a85f_b911_d7f6_1aea_1f12_2596;

        #200;
        key = 128'h014d_6cab_a54b_36ce_d9e3_d5a3_c355_a32b;
        state = 128'h4ed3_aa82_6898_557f_938c_a931_6ce9_1cd6;

        #200;
        key = 128'hba4b_7fee_a0a0_113c_8414_f5a5_d460_c232;
        state = 128'hef2c_ef80_525d_ae61_1927_0265_b287_560f;

        #200;
        key = 128'h1959_3939_6564_a46c_f620_3a25_d305_6eb6;
        state = 128'ha41b_c00d_5934_ba7d_7205_1b96_f2c4_ffb9;

        #200;
        key = 128'hfe96_7197_ced4_c3b5_6279_dda3_c90a_881c;
        state = 128'h0331_30bf_ae55_2e41_8660_498d_a7dc_cc3a;

        #200;
        key = 128'h4fc0_9129_3c52_8dd8_1dea_7578_7182_764e;
        state = 128'h4e0d_48bb_d8e2_8fc3_ac4c_412e_3200_96c7;

        #200;
        key = 128'h3fbe_8845_5d67_16f1_7dd6_16cd_d39c_c860;
        state = 128'h35d7_42e6_260a_1718_37bf_3698_0ae6_b50b;

        #200;
        key = 128'h60d2_dfed_a6cc_20f5_ee3b_8383_0565_f2b6;
        state = 128'h086f_a9aa_fa61_6121_bf5a_21e3_3e33_42a3;

        #200;
        key = 128'h873b_5a47_b8c4_4ff4_aee4_d8e8_045b_f015;
        state = 128'he9b4_810b_2042_cd1b_1677_82ab_9fdd_c2bc;

        #200;
        key = 128'h650e_5fa5_960d_eb74_55c8_c1de_c19c_c61a;
        state = 128'h25fa_9a47_1e39_81e9_9b26_c82a_72dd_a54f;

        #200;
        key = 128'h684c_0101_5e03_267c_a852_bd6d_dd3a_432a;
        state = 128'h6d12_57e1_6a0d_50ac_3ca0_6c21_99e4_17fe;

        #200;
        key = 128'h1a90_23b0_abb9_bca6_ced6_e5ef_dbc3_3015;
        state = 128'hf6a8_ab01_de66_a3a9_030e_17a5_237a_171c;

        #200;
        key = 128'hf1af_2087_e035_955d_1ee4_ba82_5f8f_eaeb;
        state = 128'h2f7a_376e_6625_7fb4_a719_7374_f9c3_763f;

        #200;
        key = 128'hf1c7_6349_ba1a_a71a_b6ae_4d7b_b031_3184;
        state = 128'h3167_30f0_91ad_b440_e3ba_cc99_2c35_f946;

        #200;
        key = 128'h7945_a8de_b72d_92d7_bb8f_6df9_90fe_37e0;
        state = 128'h150b_49f7_87cb_7d29_720c_726f_a39f_13e6;

        #200;
        key = 128'h511a_ecec_f07a_eb34_5930_a5d5_6867_e7d6;
        state = 128'h1c87_f40a_3cbf_2a54_030a_d144_b8b8_2f92;

        #200;
        key = 128'hb2e0_1795_b1de_7cb9_7f49_fbac_dd33_e645;
        state = 128'h1fea_d30b_4e12_b365_56a6_6b6f_c58e_8e49;

        #200;
        key = 128'h89da_b54f_4a10_fa6f_b354_bc56_945a_d48d;
        state = 128'hd5a9_4c15_4afa_3615_3054_a85d_e512_9c92;

        #200;
        key = 128'h7ef5_4826_8e77_119b_c0df_edd6_c90e_249a;
        state = 128'h480a_4894_ac6d_2941_2bb7_0ef1_2333_1822;

        #200;
        key = 128'hd10d_ff41_0a4d_ce4b_64eb_0436_5bc3_6495;
        state = 128'he178_80b8_8b1f_59bb_707f_05ca_3480_5d92;

        #200;
        key = 128'h2181_655b_5b87_8d2e_26b1_cc12_14a1_5a1b;
        state = 128'h2586_7401_dd94_4009_b7d4_bb29_85f2_39ad;

        #200;
        key = 128'he94c_4911_6088_eb00_ef76_6d5e_e0f1_f3f3;
        state = 128'h43ed_20b3_db6b_56bf_a477_4e72_575e_2ee9;

        #200;
        key = 128'h4c8d_5645_f177_e0f0_39d0_17f4_965a_ce91;
        state = 128'hdd30_bbc1_bc9e_b04a_5ac7_e4f8_6307_aefe;

        #200;
        key = 128'ha1f8_59b6_a829_bd39_60cd_0f77_6aa1_bcae;
        state = 128'h6b0d_d363_ecfa_0b81_d663_d1f3_07e1_a111;

        #200;
        key = 128'hbef0_03e2_a04b_8557_13c4_0a10_f3f0_80aa;
        state = 128'heca2_5712_0980_0c92_a7f0_58fc_944d_e34f;

        #200;
        key = 128'h0550_9e6d_333b_0374_f0d7_c555_92c1_4ef9;
        state = 128'h4e60_c47e_b2bf_53d9_c555_49da_9166_462c;

        #200;
        key = 128'hf97f_85ad_e7b6_0600_cf31_835c_a509_da27;
        state = 128'h6041_b22b_2239_e533_87b4_3e5e_f414_f8b1;

        #200;
        key = 128'hb7fe_c15c_af5c_e782_cd8f_5486_e7c4_061d;
        state = 128'hb965_4fcc_337a_6286_e0ae_b9fc_46f5_2e6b;

        #200;
        key = 128'h58d6_0a8c_be25_d0f5_22e1_8c85_dffd_850e;
        state = 128'h374e_32c1_dfb0_0985_3861_de9c_7547_c532;

        #200;
        key = 128'hf6ee_431a_9f5e_e247_9285_e6cf_8624_67e5;
        state = 128'h8375_f02e_5f49_3659_0748_3553_4305_2c55;

        #200;
        key = 128'hffc4_4e5b_9d0a_55b9_75fe_480b_7ec7_4e29;
        state = 128'h703f_caba_32e7_157c_3daf_320d_e842_587c;

        #200;
        key = 128'hf7a1_9162_671f_0778_7b12_5042_e1df_c36c;
        state = 128'h3ea1_fcd1_8eb6_da08_d581_54eb_c117_649f;

        #200;
        key = 128'h1b5a_b871_62b5_9902_ab74_10bb_53ed_1b9e;
        state = 128'h7c23_e954_3811_ad58_29ea_09d8_7a68_61ef;

        #200;
        key = 128'h0030_541c_159a_ec61_f8bd_6beb_7670_a1d0;
        state = 128'hcb9d_9586_3f8d_9dc8_c900_1271_1caf_6b69;

        #200;
        key = 128'h1fca_e96a_8ed9_c6bc_6b90_5557_11ce_63b7;
        state = 128'hbafa_4269_8ddd_6d45_6ef0_223f_fcad_ced1;

        #200;
        key = 128'h6cce_232f_bb3f_9dea_16fa_f852_7954_739a;
        state = 128'h26ec_682f_91b9_bc6a_7035_5ce2_0e19_0772;

        #200;
        key = 128'he6fe_f39b_407a_9af6_a952_3c99_e71f_f19a;
        state = 128'hfe53_3209_6a03_8ce2_e4c8_b706_7156_210a;

        #200;
        key = 128'h931d_e8c8_fa6d_5a58_a655_d4f1_4ce5_a143;
        state = 128'hb5ce_a9b4_b4cd_048a_2d4c_7658_2d01_b3c8;

        #200;
        key = 128'h6623_9442_2186_b91e_78ba_8cb8_90ef_08ce;
        state = 128'h9518_1a10_6c25_a6fc_1e03_00af_5ecb_4e0b;

        #200;
        key = 128'he39d_9afa_e0be_8bb0_c607_3d34_4eb1_81ac;
        state = 128'h2065_8e98_0cbe_f289_8a89_75cf_499f_117e;

        #200;
        key = 128'h887b_0692_3416_90ce_61e3_1e77_4279_eea4;
        state = 128'h9e8f_57c8_6417_146c_ba87_f5e0_50fd_d5fa;

        #200;
        key = 128'hb0ee_d887_7407_39b7_e2fe_2dfb_f226_4701;
        state = 128'h3832_a410_e18f_0f1c_cc5a_057a_efb1_6bab;

        #200;
        key = 128'h3a0f_f405_71b1_ec36_fa53_1ed3_9041_e1e3;
        state = 128'ha0ff_3a23_0656_02f1_40e6_6ca7_8e15_977d;

        #200;
        key = 128'h19b4_a5c7_d5d9_2e32_47a8_11c6_9b93_f30e;
        state = 128'h6725_92e3_bfae_c2a9_951e_22ae_74ec_a764;

        #200;
        key = 128'hf7d6_f2e2_134e_aff2_43e2_2c51_9ada_3f06;
        state = 128'h1531_f924_9dfc_a8b0_6591_9d2b_85fb_4fb8;

        #200;
        key = 128'hb16e_74ba_9217_d24b_72c8_5651_fde4_f4d1;
        state = 128'hddbe_4cab_0825_e32a_0da7_6da7_9a24_bebf;

        #200;
        key = 128'h9776_1c6f_3ebe_c87d_a137_35b2_5b35_cc2b;
        state = 128'hd7c4_41d2_1f63_54ca_6edd_18dd_fe41_736b;

        #200;
        key = 128'h56ec_34ca_d8bf_6c4a_5643_e901_0d26_8d75;
        state = 128'h2830_d167_372e_7c65_ce40_78ec_a834_f07c;

        #200;
        key = 128'h35c3_be20_0eda_2993_4bc4_d099_8f9a_1a3d;
        state = 128'hfafe_f2ac_0b84_aee9_8da2_2787_c4db_e0f8;

        #200;
        key = 128'hb3c1_b532_d065_7a9f_faf1_f145_6e30_db9b;
        state = 128'h351e_fc85_a257_8c3b_89e5_158a_9838_3af6;

        #200;
        key = 128'hf6b0_29de_58fe_fd5a_a509_6148_ef88_11ad;
        state = 128'hd5b4_5ff6_5236_7ba8_1fc8_e1ad_bfa7_b3e0;

        #200;
        key = 128'h1081_3cd3_8df0_f55b_27d4_31e8_4a96_1b45;
        state = 128'hcca2_fbd1_42e0_c567_02d1_66bf_2d7c_688f;

        #200;
        key = 128'h4dc8_51ca_e1a7_4d0d_d372_d3fe_8cf6_9e71;
        state = 128'he59a_78c0_1822_1ebb_7a88_5b9a_a1dc_fd96;

        #200;
        key = 128'h694d_192e_a582_f27f_ef34_b8d1_4024_2f06;
        state = 128'hcd90_1463_c40e_f88a_498e_dc01_1ae3_5a61;

        #200;
        key = 128'hcf4a_4387_4c8c_6266_27f2_7c91_a6b8_0d69;
        state = 128'hb876_f56d_c711_cb57_a009_47a4_43c9_06a6;

        #200;
        key = 128'h63f1_f126_4271_2460_855f_db9d_f193_988e;
        state = 128'h86e3_bcbf_7493_4531_5cdc_37cf_f1d1_7cf6;

        #200;
        key = 128'h58e4_30b5_87a5_082d_8edc_6487_ebab_30dc;
        state = 128'h6d2d_91fa_35f3_bc28_06a8_106a_bcf2_63ce;

        #200;
        key = 128'h22b6_1884_d83c_35d4_6749_558f_a7fc_2f4e;
        state = 128'hf0c6_8dcf_9a1a_5f42_7984_3494_95c4_8d1d;

        #200;
        key = 128'h46ba_01f2_ee09_4300_57db_7859_b817_1e77;
        state = 128'hbbe7_478e_31b0_8110_92b0_5eff_ea59_6c5e;

        #200;
        key = 128'hd078_341a_f2cc_565f_98db_279d_0f66_21fa;
        state = 128'h0749_7c72_7691_a92b_b133_9468_918e_4c70;

        #200;
        key = 128'h2ad4_259e_1089_ab5f_97fc_a2a9_eb44_0f5d;
        state = 128'h3c75_a5d8_07fb_ece3_20cb_2976_1f4a_c0e6;

        #200;
        key = 128'hd114_bcb5_a9e3_fc27_5cc0_efa0_cdd1_2b93;
        state = 128'hf4fb_8694_1250_3aad_6928_f1c3_d40f_1182;

        #200;
        key = 128'h5418_cb30_2543_5eae_47aa_5214_58b9_cd2c;
        state = 128'hc3e2_0913_c026_e939_bf94_15a7_f183_63d7;

        #200;
        key = 128'h9b60_8c93_b5a3_c9c3_e2bc_f38a_2977_0e6c;
        state = 128'h4c10_c3fc_237f_212f_1c1f_0ddf_87ce_34d5;

        #200;
        key = 128'ha01f_a350_a150_3015_d8dd_d943_bded_7cac;
        state = 128'h03c5_705f_98f7_ccfa_8673_5750_8990_0e87;

        #200;
        key = 128'h7f0f_5126_eed2_b7a1_aff6_db8c_3659_34f6;
        state = 128'hf2f2_565b_7b29_e2e8_b2e7_0209_b28a_f09c;

        #200;
        key = 128'hba80_183d_8b3d_4949_76a2_6286_71dd_494d;
        state = 128'h7385_bab7_6cb4_e75c_70cb_3c3b_77b3_6ba6;

        #200;
        key = 128'h2c5f_4ffc_dad5_d6d1_9521_e7fe_eafb_c10c;
        state = 128'h634c_243f_101c_0070_e8e4_3dc9_874f_ddac;

        #200;
        key = 128'h761b_07cc_135f_1313_0676_683f_5e86_d84d;
        state = 128'hcb13_d392_838c_b22b_c983_0bd7_a072_e831;

        #200;
        key = 128'h8abd_503b_f79e_8b28_5d91_8e5d_0b01_3bb5;
        state = 128'ha197_1087_3562_c7d4_5890_5f2a_494b_408a;

        #200;
        key = 128'h8c17_9864_5d51_278a_6435_61d1_7398_15c7;
        state = 128'hadd6_d0c7_128b_c3cc_1d1e_8e51_f841_6b76;

        #200;
        key = 128'hf9c9_81d8_9bf7_a802_3319_e442_8e1a_42b6;
        state = 128'hf417_015b_a3bb_2f2b_27ef_1643_6ddb_f27a;

        #200;
        key = 128'hb250_b6e2_c09f_745b_8121_d794_558e_f019;
        state = 128'h6531_b281_5adc_8a7d_78a1_84c3_3469_8f0f;

        #200;
        key = 128'hb1e3_21e3_e83c_c58c_7609_7089_0220_845f;
        state = 128'hab43_2fd6_2019_ba4c_3a42_a8c0_bcaf_cba2;

        #200;
        key = 128'he85e_2497_1a0a_f1f4_26f6_f554_aa6c_3a18;
        state = 128'h10d4_f3a7_1ca0_791c_c2d2_ff40_e851_fb51;

        #200;
        key = 128'hc686_ac53_aa2a_8bdb_21af_c583_8f93_b58c;
        state = 128'h968b_3ac5_8c08_8d9b_3e88_3889_b1f3_242f;

        #200;
        key = 128'hfa8a_dd93_f398_59bc_ddca_724b_12e2_aa3f;
        state = 128'hccbb_4bde_8f29_fe3b_4fe1_0acd_25c5_5f53;

        #200;
        key = 128'hf1b4_0dfc_2b02_bad1_f0a5_2e57_d718_7491;
        state = 128'he47c_81e5_cdd4_c6a7_b2fc_493e_98f3_3246;

        #200;
        key = 128'h71bf_b262_c308_19e2_3b09_5170_e25f_fd73;
        state = 128'h373f_f48d_257c_454b_915a_e9f3_f083_7109;

        #200;
        key = 128'hb050_69f4_5b5e_a68d_a61c_82de_9324_0439;
        state = 128'h1163_996f_16f2_f05e_ac6c_78dd_1573_1eb1;

        #200;
        key = 128'h414a_fb21_a92b_464e_b5c6_fbd5_9bf6_2ce7;
        state = 128'h90b5_f517_24f4_3cef_1675_669f_7f41_9380;

        #200;
        key = 128'h2441_8526_9bb3_ffcc_dcc8_b807_e012_c2dc;
        state = 128'h161d_5f2f_7f37_b0bb_41dd_4578_8fc7_e6db;

        #200;
        key = 128'hab84_8f6b_995d_a696_b6e5_b1b2_30b9_1c15;
        state = 128'h7e6d_3c08_674f_aa43_7fdc_40c8_7845_72d9;

        #200;
        key = 128'h4e9f_76cf_0ed9_a69d_c00c_f343_77bf_1310;
        state = 128'hb476_3fff_36fe_1e05_d64b_56d2_3c16_a236;

        #200;
        key = 128'hce26_200a_4853_390c_8b48_05d3_4a25_8fd1;
        state = 128'h5445_e9b0_a28d_cc84_eaa8_e934_6ec7_a6f9;

        #200;
        key = 128'h3fd7_d5c2_36dc_68bb_33da_ebfe_566b_3430;
        state = 128'h1d08_54d6_1e4e_01ce_5f78_d044_75ff_d4b2;

        #200;
        key = 128'ha55f_2dd5_7f5e_3922_dd79_33b9_872a_795d;
        state = 128'h82b4_c64e_4308_b0a0_c811_d726_ff67_bb59;

        #200;
        key = 128'h13c9_f346_23fa_f26e_5c2b_0ac3_d843_e46b;
        state = 128'h08f0_f243_17d7_14cb_b1f7_b0d8_a573_3eb6;

        #200;
        key = 128'hac20_2bac_8e94_f302_6c8e_400a_fc66_94f2;
        state = 128'h4bcc_eb26_b200_1542_5559_9003_fb82_5064;

        #200;
        key = 128'hf369_3cd3_d53c_f37a_1fc9_0335_79a2_28ef;
        state = 128'h196a_1c54_19df_df56_3be1_69be_7638_7d72;

        #200;
        key = 128'h059b_65ad_6813_e4a2_7d1c_677e_2d68_c95f;
        state = 128'h2877_cdd5_df3f_87b1_ae55_a348_0227_32fa;

        #200;
        key = 128'h443a_6895_791c_aa12_25f6_d78f_1d8e_3e80;
        state = 128'h5b60_3a2c_c50c_d807_3a7f_12b7_69e3_9601;

        #200;
        key = 128'hb4f2_bdb1_ba80_8d7e_b335_3a9b_8a6a_2eb8;
        state = 128'h3611_a122_50ff_f53c_a0a6_4f0b_3518_00a2;

        #200;
        key = 128'h0eb5_aa8c_029d_66c6_585b_0b35_14ad_bcad;
        state = 128'h4c31_5000_e9f9_9dbb_1df8_1297_1e22_e8be;

        #200;
        key = 128'h4ae3_8f00_d38b_a008_f785_0769_2696_17fc;
        state = 128'h02a3_2199_0d52_8109_28a6_be42_feba_f0f5;

        #200;
        key = 128'h9ebb_6d83_4c1c_46c8_5f58_b4f9_8c3c_a454;
        state = 128'h411a_c4a6_bbee_1b9a_8d28_dc2d_00fd_140d;

        #200;
        key = 128'hc934_e2da_3166_d8f6_56c9_197c_602c_7c73;
        state = 128'h58a4_0e3f_eeec_3478_7915_19bc_149b_2efd;

        #200;
        key = 128'h7243_e2d9_b710_f702_c903_28a7_04ed_1c1c;
        state = 128'h06ee_f71d_60a7_1d65_b347_5c9f_1893_8fd4;

        #200;
        key = 128'hac7f_2c74_d790_9eef_b27c_0ea8_b25b_bcd8;
        state = 128'h9fea_bef9_3330_d241_100b_dc1a_0db2_4b3b;

        #200;
        key = 128'h6b20_202b_f5ac_1d23_0a36_26b2_3f51_4398;
        state = 128'h78e6_d0b9_d7cf_f258_b2e6_ea14_dc09_5a84;

        #200;
        key = 128'hdead_693f_a2cd_f028_f106_be4b_93f4_d285;
        state = 128'h2b27_719e_8aa4_5137_ffaa_e42f_26ba_4832;

        #200;
        key = 128'h6fcd_57ba_2dcb_21e1_cce4_2bb3_e4ef_4dce;
        state = 128'had05_1590_d4b0_64b2_30f0_87d3_d63f_685c;

        #200;
        key = 128'hb5be_d067_fe23_9295_7b4b_d14a_ec20_6090;
        state = 128'h12c2_bb7d_fae8_3caf_795a_9c61_a1f3_815c;

        #200;
        key = 128'h9d1d_c99f_67f1_da57_13fa_1c67_b1ae_d20c;
        state = 128'hfc71_a470_911b_38ea_91e7_ef8b_ee3d_a93c;

        #200;
        key = 128'h3ffc_1aae_754b_0853_774b_d373_d41f_efec;
        state = 128'h5daa_8894_c96f_9a79_0c3c_5652_6c96_9da6;

        #200;
        key = 128'heaaf_407a_6db9_a6ce_b2ea_efe7_fda2_3c50;
        state = 128'hd9c4_3a34_deaf_9966_2c8e_f2f9_c91d_2d4c;

        #200;
        key = 128'h46e8_b92f_6b25_b8a8_6e18_a134_9039_e673;
        state = 128'h0ccd_3252_792f_c301_b0c7_d903_a795_dcb1;

        #200;
        key = 128'h3257_d9af_624b_ac47_5f7b_f446_f5c6_c869;
        state = 128'hc2c6_39b9_c111_b802_d53b_70df_4876_115d;

        #200;
        key = 128'ha782_c9a5_383f_1055_cb62_147d_858c_3fc4;
        state = 128'h12e8_19b6_a2d7_36e2_8394_49ff_0c77_7f04;

        #200;
        key = 128'h1183_770e_32f8_6a8b_c89e_4af3_5beb_02c0;
        state = 128'hc2e4_b6af_3ff4_e9f0_6c94_5566_47af_8ffd;

        #200;
        key = 128'h4187_423a_7398_ceae_2f53_4b87_a582_f413;
        state = 128'h7414_1300_7eb4_bac0_013c_6ebe_d325_3e76;

        #200;
        key = 128'h43c1_a93a_a16d_bd08_6637_69ab_da35_d51f;
        state = 128'h9568_9deb_b0f7_3b08_9b80_7db1_1236_1eb0;

        #200;
        key = 128'h7a9f_0a11_a471_b0dc_a7e1_6118_1d43_366d;
        state = 128'h9d99_bdec_daa6_a1df_71b6_1a15_08e9_fe79;

        #200;
        key = 128'h8b84_3681_bf2c_7384_574f_37c1_000a_c083;
        state = 128'h368f_5cb2_4837_6922_7ce4_d6e9_7b2d_0d93;

        #200;
        key = 128'h0a21_b9fb_bbf2_4336_e54b_ffd9_0751_f3bf;
        state = 128'h1409_01ce_7247_a3fe_c01f_d391_2f69_a039;

        #200;
        key = 128'h4226_7015_2f42_db9b_ec14_4c5b_8cdf_8f41;
        state = 128'h38a5_4ea5_0c7a_600d_0e98_90dd_da62_ed5d;

        #200;
        key = 128'h83a3_3b7a_8ab0_579b_9eba_8ee2_0e06_e4b8;
        state = 128'h901f_d4bd_998a_3a02_a5d4_e139_5c0f_5645;

        #200;
        key = 128'hdab1_5b36_61cd_0598_3a39_9f82_0b08_ff9c;
        state = 128'h0776_6e53_f9a2_0efd_56ac_7c04_7553_0f14;

        #200;
        key = 128'hae0c_03ba_d1e2_707d_23b0_d78a_273a_fa9c;
        state = 128'h5183_c8cb_1089_c16c_eaf2_73c6_afc7_4984;

        #200;
        key = 128'h6cdd_9694_976e_36bd_02d0_3e82_49fd_e2fb;
        state = 128'h01af_2944_6232_9182_28af_1751_83d6_211c;

        #200;
        key = 128'hc8e0_d10c_5652_529d_a72e_a006_750d_7dfc;
        state = 128'hbee4_bb12_d827_807c_b109_bc5c_ec10_bb7d;

        #200;
        key = 128'h4c33_9ea7_f14f_db51_93ad_41ef_9da3_2692;
        state = 128'h1307_ea4f_f2f5_43e4_7d07_e3e5_1bae_1b0f;

        #200;
        key = 128'h10f5_0a13_6c39_c9a7_937b_4dcb_03cc_1546;
        state = 128'h9c5a_ae8d_d48f_7ec8_f40b_9fcf_92de_69bf;

        #200;
        key = 128'h1d48_cfd3_bafd_8fe8_7b01_dc8c_a39d_f88a;
        state = 128'h8f09_99ca_f589_c2b7_23e6_28e8_6a6b_568f;

        #200;
        key = 128'hfb72_ee43_d5ee_cede_cb71_e01a_1b50_0471;
        state = 128'h37e2_d7af_3dae_f890_172f_b0a0_7a69_3f63;

        #200;
        key = 128'h6a83_5878_64b7_a681_725c_ba91_ca8a_9598;
        state = 128'h9ed0_34c7_96e5_f7b8_0b4f_d042_c29b_b43d;

        #200;
        key = 128'h6fda_d13b_01e4_43c4_209e_d4fe_2571_6424;
        state = 128'h2316_1f6e_443d_a963_3437_d673_c996_483e;

        #200;
        key = 128'h28d6_1a05_7100_3b04_16e3_a447_3cca_f0c7;
        state = 128'h5aec_56b7_d57b_5777_c98d_a40d_a56a_95d3;

        #200;
        key = 128'h0d8c_9c64_eb39_c614_52b7_2483_fbbc_66d0;
        state = 128'h1aee_91b9_e0a2_622e_24b5_3bdd_c5b3_54b2;

        #200;
        key = 128'hd3f3_6ba4_d110_69dc_6b19_05e0_946c_c120;
        state = 128'h98de_dd55_9abb_4779_d3db_30cd_546a_4b46;

        #200;
        key = 128'hcb9c_361d_bc96_c15b_b4c1_c560_54d6_fbaa;
        state = 128'h6a6f_8201_2247_7837_26bc_6472_2592_fa24;

        #200;
        key = 128'h3660_e8b4_6131_f93c_8e38_05a9_46e6_0e7b;
        state = 128'h5df3_925a_315b_d53b_882c_6030_0e1f_4815;

        #200;
        key = 128'h3140_a99c_3012_64f1_2ed5_df47_69e8_c100;
        state = 128'h3375_241b_ccfb_9614_322a_a508_29c7_38ab;

        #200;
        key = 128'hc1be_7705_82ae_5230_38a4_380b_2a1d_4d8a;
        state = 128'he328_2b82_afc7_2bfd_39f7_9674_c899_c2b7;

        #200;
        key = 128'h8bae_6b91_997f_8732_c4bb_aa35_5a82_9125;
        state = 128'habe6_7c6f_87da_c512_7b3e_6700_7bbb_d050;

        #200;
        key = 128'h0ee4_cac4_0d30_3790_9617_bb10_f683_a65c;
        state = 128'h2d88_573a_bb82_753c_7aa9_091e_6a56_de83;

        #200;
        key = 128'h1f29_1ac4_b25d_7ae6_ba05_984a_db87_a06f;
        state = 128'h4b01_28b8_f336_fd30_b9ac_31a3_c86a_b782;

        #200;
        key = 128'haca8_6792_2aa5_73cc_8ead_c0c7_508d_a1bd;
        state = 128'h5e0b_5478_e2b4_01bc_300b_7bb3_32ae_9334;

        #200;
        key = 128'haceb_6b29_0a8c_ec93_6c50_55a8_6ec4_edec;
        state = 128'he797_f09f_266e_96a5_22af_510f_b69d_c495;

        #200;
        key = 128'he7b1_9fe1_3427_9dc1_01b8_3333_6bd5_6339;
        state = 128'h94d0_b2a6_64e8_36c4_7fde_4cb3_edd2_4604;

        #200;
        key = 128'h89fe_0b27_ddd8_86ae_a0b1_2ffb_c1b7_689b;
        state = 128'hbc15_9fe5_cac0_3ef1_516b_5d97_7d7f_bed9;

        #200;
        key = 128'h13c1_4020_efa5_bd86_d7f3_badf_aafb_4f6f;
        state = 128'headd_a481_6bff_7600_0d15_ed95_f8b6_6625;

        #200;
        key = 128'hd185_766e_5488_30ad_2052_4561_b775_d6de;
        state = 128'h9901_63a1_00d5_70da_b5b7_80a8_7f64_aa64;

        #200;
        key = 128'h1c2c_4e54_ff37_874b_8093_dfea_6340_3095;
        state = 128'h2771_c08f_99a7_3409_57d4_db9f_627d_24df;

        #200;
        key = 128'ha13e_4193_6be5_dca8_5945_469a_f3e3_4621;
        state = 128'h9cae_6397_663d_5f45_e7df_2098_cf52_1ccd;

        #200;
        key = 128'h4086_81e4_c293_6719_f3fe_5e9c_8615_bda6;
        state = 128'h5608_ee0a_c9a4_8d2c_f835_1a02_f437_2135;

        #200;
        key = 128'h6ff1_17c7_ac1c_47d5_5c68_34b0_e4c2_9349;
        state = 128'h9beb_3c0b_de1c_841c_1ab1_f5ef_0a75_1868;

        #200;
        key = 128'hf582_25b5_c1f1_87cb_324f_8972_4bec_e76c;
        state = 128'h9947_bb15_06c0_9bed_97d2_de94_e156_a86b;

        #200;
        key = 128'h7e17_c286_f9b6_8624_60c3_1df2_19c8_14b5;
        state = 128'h7c9f_2617_34c2_23de_3f2a_f819_a8c4_7563;

        #200;
        key = 128'hfa30_472f_a20c_164f_464b_3610_f92b_10bf;
        state = 128'ha31d_c194_2130_e6c2_33b1_62be_7605_a51f;

        #200;
        key = 128'h345f_d59b_0365_1bac_b6de_cc6a_e5d0_56c0;
        state = 128'h37cc_b860_49c3_0f27_a036_d508_4831_c6e4;

        #200;
        key = 128'h7b9b_af2c_15f6_45f1_7807_c746_0e64_2048;
        state = 128'hd04d_2547_5428_859c_7efd_e955_f693_f6f3;

        #200;
        key = 128'h56ce_8e6e_316d_2c89_6929_6c5a_fe0e_f08f;
        state = 128'h25a9_fe8d_c653_5e2e_7541_f01d_145c_8657;

        #200;
        key = 128'h681a_8de2_9a8d_f7fb_1564_bf28_fbcd_6a5d;
        state = 128'hf156_0445_8795_a287_6672_ae3c_a1d5_2158;

        #200;
        key = 128'h980d_4742_7d76_2fdf_f0d7_71e8_1202_5d32;
        state = 128'he21c_f342_d11a_37a3_5dd7_d22f_8216_01ad;

        #200;
        key = 128'hf125_8559_bf18_5ebe_87f4_8416_5b22_a882;
        state = 128'h8327_9d23_5b8f_2888_746a_40b9_f5dc_74c7;

        #200;
        key = 128'hf6d8_fc4c_4ea0_9e4f_3594_f98c_9211_dd97;
        state = 128'h3523_fe00_4115_87e0_8024_05b8_ec19_8ca0;

        #200;
        key = 128'h037e_a96f_0672_9328_c5c4_c54e_8fe9_a2e9;
        state = 128'h67eb_30ff_af20_48c1_4cf7_e9d8_25dc_eb63;

        #200;
        key = 128'hc772_da88_fc6f_9615_4247_1928_8ef7_9003;
        state = 128'h2b9b_2eaf_9d9b_3393_48d0_9f8f_2edf_68a5;

        #200;
        key = 128'hcec6_80c7_c3c8_b3f6_aa1b_2022_b2b3_8e8c;
        state = 128'he116_7ad3_b0cc_b13d_05e5_4d90_bdd9_4af8;

        #200;
        key = 128'h765a_ac34_910e_ce96_6f79_c062_1d56_3454;
        state = 128'hc0ec_90aa_84cc_209e_14a1_7e10_dc36_0d60;

        #200;
        key = 128'h916b_c4a2_b968_ee49_bfd1_b61b_6858_72e4;
        state = 128'hdbf9_dd06_91c2_efa2_6bc9_11d1_d05e_7d85;

        #200;
        key = 128'h9aa7_2102_fd11_5d6b_1bc1_08e9_2278_281a;
        state = 128'h5a3c_a6e3_e937_bbe9_0fcc_f0a8_e55a_0c33;

        #200;
        key = 128'h21d2_865d_b498_5625_a479_2439_992a_a793;
        state = 128'h4acb_2203_95c6_6928_ab29_373f_b071_3e42;

        #200;
        key = 128'h84b3_75f7_1a81_33f3_d749_801f_9310_4640;
        state = 128'ha994_f091_1887_3c3f_4c78_9893_33ff_7cbb;

        #200;
        key = 128'h0050_5772_6f34_480f_70da_3e39_15a2_e53a;
        state = 128'he90d_a80e_9af9_f570_82f2_5ff8_d7c8_588e;

        #200;
        key = 128'h21ff_e991_5edb_14f1_2b2d_fee3_5657_dbfb;
        state = 128'h6c2c_3747_476f_7437_a77f_6eef_0d6e_b375;

        #200;
        key = 128'h7c11_d84a_8449_c26d_48bb_390d_ed1b_234b;
        state = 128'he34d_f78b_352f_aca4_f026_de0a_4cee_7f0e;

        #200;
        key = 128'ha129_e49b_1e04_03f3_40d9_f81c_ec19_f437;
        state = 128'h5104_ee22_54ac_0ea0_d12d_134f_e980_a2ab;

        #200;
        key = 128'h28f7_614d_0090_92dd_9142_a956_a29c_0b27;
        state = 128'hfc71_319f_9195_c569_c718_187d_84cb_da8b;

        #200;
        key = 128'h12ad_4687_33cb_0258_9c2e_8391_ce10_93e8;
        state = 128'h6f8e_190a_968a_daaa_e820_9535_c263_610a;

        #200;
        key = 128'h73d2_e2b5_5b61_fbaa_f7c4_9a1f_2b39_04cc;
        state = 128'h03bb_6b9d_71b7_3591_61bc_6f4e_28d3_3aae;

        #200;
        key = 128'h7f6d_8c53_fb6a_47e9_b15a_02bf_c353_7cdf;
        state = 128'hd044_0252_abb1_470b_c723_07a5_ef57_7029;

        #200;
        key = 128'hf60f_7ce0_34d2_2105_2683_0eb7_caa8_1622;
        state = 128'h0f4d_6254_bc43_5037_a796_a799_9e0d_060b;

        #200;
        key = 128'h46ac_11b8_9c03_310c_f67d_6a5b_0f7f_f95a;
        state = 128'h59c6_46a3_5d2c_74fe_c049_8d89_bc1f_4822;

        #200;
        key = 128'h693c_0683_e43b_3f38_e7ff_cd93_f340_9676;
        state = 128'h07dc_9aa2_5f75_8e85_f179_b240_1474_2632;

        #200;
        key = 128'hdeb3_7bed_ee5a_5b01_2249_b615_192c_7f6b;
        state = 128'h67af_d526_5452_1d56_84e8_efb1_c587_2fd6;

        #200;
        key = 128'h84ad_f765_5016_7d15_b3e6_9968_7d9a_9e02;
        state = 128'h3649_2ed1_0a2a_ed4c_c065_fc35_f22a_d8f6;

        #200;
        key = 128'h0fb3_3f74_47cc_4a38_b000_4d8c_189c_d4f9;
        state = 128'h7746_37d5_3ee3_0d5b_9111_7740_7bd1_4537;

        #200;
        key = 128'hc0c0_55f9_5bdf_76b2_55b2_5751_b2ea_40cb;
        state = 128'h3a8c_c61c_0550_9f0d_0e5a_dc5a_ec62_35dd;

        #200;
        key = 128'h122b_b505_0733_fa52_8c36_18ed_2a71_c8a6;
        state = 128'h2f95_5c60_d96e_e6ec_865c_1f3f_ab5c_70dc;

        #200;
        key = 128'h5a3a_d3ce_bae0_6f02_d8ca_94d3_9d92_6700;
        state = 128'hbfd9_18b2_4251_3298_83ed_aeb9_41c1_538a;

        #200;
        key = 128'h7453_6a78_cb4b_1089_f504_f181_afdb_4b64;
        state = 128'h474e_1181_bcf9_bcae_08b6_7545_47f2_0bc2;

        #200;
        key = 128'ha5b6_ffed_8d10_222e_89da_ecfe_783d_2f0a;
        state = 128'hc934_aa1b_3cd7_8953_dac7_4b1a_48a2_8c36;

        #200;
        key = 128'h26ac_ce25_c5ed_4bcd_6c2f_4aae_c08f_d544;
        state = 128'h5ff5_9794_6112_2c32_f09f_45a6_825f_4b0f;

        #200;
        key = 128'hf0f2_13af_a827_a17d_eb17_7081_0e4c_e054;
        state = 128'h6202_3625_94f1_d6e9_5ed0_281d_ae9b_1797;

        #200;
        key = 128'h0af0_a986_3569_18f0_f418_7256_b570_5dd8;
        state = 128'h14bf_5cad_4b79_5f67_a976_eebe_702f_720a;

        #200;
        key = 128'h22b5_7c55_c74f_47d1_541e_717b_84e9_6f0b;
        state = 128'h9cdc_f431_5253_2dcc_3b90_974e_5258_f62a;

        #200;
        key = 128'h53c7_0162_b93c_d3f2_7f18_0768_cf64_9893;
        state = 128'h7504_6f0f_61a7_70fd_607d_5996_cccb_8910;

        #200;
        key = 128'h1014_5ffd_96ab_7875_dcb5_4349_6a6a_11fc;
        state = 128'hbfce_db00_e853_c41a_a280_192b_ac7d_b664;

        #200;
        key = 128'h502f_b8dd_be2f_c667_32e0_c8f9_14f6_88de;
        state = 128'hcfa9_78e0_dbed_7353_d78a_cfd0_e706_1d7b;

        #200;
        key = 128'hf12d_c72c_1abe_246e_6ffd_ff16_3c0c_a4a9;
        state = 128'h54b9_5a7c_3343_7060_fdf9_b5f0_86b7_9e95;

        #200;
        key = 128'h4efb_202e_5433_6dfa_0518_81af_5934_d721;
        state = 128'he9f9_dc04_204b_c5ba_cfe1_12eb_d2de_e044;

        #200;
        key = 128'h72f3_7327_19bb_137a_2131_f756_0423_53f9;
        state = 128'he63a_f298_5bf0_d111_4b4e_0a33_99d9_07e0;

        #200;
        key = 128'h7371_478c_f2b0_3a37_3267_78e1_f99f_a3a5;
        state = 128'h3f71_69df_d55b_8d77_503f_72e4_43de_8656;

        #200;
        key = 128'h6e4a_67d8_bb6a_7d65_1d91_8dfa_dea0_08e0;
        state = 128'hca73_593c_b078_cb33_5c26_4120_a1e1_ca3b;

        #200;
        key = 128'hdc4c_4e3e_22cf_f338_db9b_715f_b18e_c919;
        state = 128'h1ab3_d4b5_903b_dd8b_9473_3438_439b_563c;

        #200;
        key = 128'he45f_d67f_5d1a_23d5_a57c_b6be_ccd9_5973;
        state = 128'h3b54_105e_33a1_7b66_591b_4a84_437c_4399;

        #200;
        key = 128'h38f3_844b_6898_3f8d_44b5_7169_42a4_1c09;
        state = 128'h2864_6a45_a9dc_0df9_3b4c_88c0_396c_5e82;

        #200;
        key = 128'had9c_04ec_0066_0c6e_a4fb_330a_fb9e_851a;
        state = 128'h5543_473f_aa5a_6d45_e559_7d3b_0e8b_bfc8;

        #200;
        key = 128'hfbb3_57cf_fdbe_e0ea_3bf5_a46d_ca1d_a31d;
        state = 128'hc7aa_a842_f1a5_71a2_7d89_816c_a7e3_f04e;

        #200;
        key = 128'h3528_037e_e0c0_e6dd_2a2a_1285_a95f_db9d;
        state = 128'hd151_67bb_e983_4f96_928b_075d_f856_d707;

        #200;
        key = 128'h2748_d850_e6fd_9c09_ebd8_f8d8_8b6b_89b7;
        state = 128'hd9cb_29e2_ba54_f787_b47f_4ee1_0cd2_1cb5;

        #200;
        key = 128'hb613_973e_60a9_9414_8070_590d_b7ac_26d6;
        state = 128'h5e52_7699_d9c6_fe9a_07ff_2ccf_beba_56e1;

        #200;
        key = 128'hc36f_59a3_58b1_e7df_8416_c874_476d_f509;
        state = 128'h5522_bebd_f7c2_d621_b570_cbf9_0a65_a6e8;

        #200;
        key = 128'hf0fc_27d2_ca90_3e53_a10a_29a9_f068_d536;
        state = 128'h22bc_a915_eced_3122_2056_b7fd_d7b6_6e66;

        #200;
        key = 128'hc057_5b91_4080_319f_290d_da7a_6228_137e;
        state = 128'h70f3_f550_9ed9_bc4a_046a_c607_cadf_a097;

        #200;
        key = 128'h1846_79c3_60a9_1adb_270f_6808_415f_033a;
        state = 128'h2db1_e0d4_128a_3b06_701a_d3ab_9e20_c3e0;

        #200;
        key = 128'h186b_515a_ca9f_6f45_4cc9_9880_151a_92bd;
        state = 128'hcea9_fa83_c995_c282_057e_324c_71b2_8296;

        #200;
        key = 128'h698f_36a1_87fe_3628_9703_b3da_37e1_56a3;
        state = 128'h9025_262c_114b_58ff_2f72_15c9_c164_fdb9;

        #200;
        key = 128'h0568_7afc_4e91_b029_cabb_237a_8ddb_eb72;
        state = 128'he2b4_c812_8f2c_ec86_d138_c539_d743_dfe7;

        #200;
        key = 128'hbed4_e288_631b_4800_fbcd_0631_6f54_c21b;
        state = 128'h7cc8_7a54_9661_3ffb_07c6_fc15_5217_4955;

        #200;
        key = 128'ha3dc_2384_2328_dad5_c718_1a27_b47d_878d;
        state = 128'h3a4d_b100_32a6_ea04_b43a_7c28_5906_70ae;

        #200;
        key = 128'h2239_1a51_7cef_2a67_b4db_e6f7_2f7b_051e;
        state = 128'hd296_abd2_da54_17a7_8013_0534_b650_1372;

        #200;
        key = 128'h2571_7cef_3d9f_6081_8d4e_bfc6_1d61_c42f;
        state = 128'hb222_89fe_9461_f831_5634_19a8_2934_f8a4;

        #200;
        key = 128'h9258_83ce_6bc3_ace5_03bc_3da3_3d50_d75d;
        state = 128'h11bf_8899_8dd1_c1df_95bc_1e74_e137_782a;

        #200;
        key = 128'h2c09_b99f_ee0a_7605_fd69_cf33_ebde_c990;
        state = 128'hc67b_917f_f162_c52c_ab98_0eff_4200_6d21;

        #200;
        key = 128'hdd9b_1a43_fec2_117e_2cdd_744c_d635_fc52;
        state = 128'hd2cc_7c52_9b4c_f711_218a_4471_0940_04bc;

        #200;
        key = 128'h11e6_8a9c_2197_0706_545d_cffb_65e6_bb2f;
        state = 128'hdb0e_7bbb_a53b_8f04_9198_d969_cd3b_b488;

        #200;
        key = 128'h9b78_3579_809b_1825_e05d_cba0_ee7b_c950;
        state = 128'h5bbb_0c72_2c10_3f80_69aa_b9c2_ded7_b532;

        #200;
        key = 128'h6754_9d96_0dd9_c6b2_0072_88cd_7466_1824;
        state = 128'h808e_e681_639e_3c4f_beee_b218_8d90_5264;

        #200;
        key = 128'h175d_6b1b_855c_a671_9d74_439d_c9d0_d461;
        state = 128'h084a_4e62_9755_21ba_c959_5e4f_c15a_e285;

        #200;
        key = 128'h4311_da4a_5ac5_d6db_5086_948b_ac3e_1ab7;
        state = 128'h33d3_8372_2d76_6409_477e_5803_8eaf_e17d;

        #200;
        key = 128'he5b2_0e68_3e7e_8b54_d36d_7bab_df80_bb76;
        state = 128'hedaf_8ea5_f092_e3f5_7140_bfc7_56e1_52ce;

        #200;
        key = 128'h6d22_dcb9_4afb_865a_4d0c_050e_7b41_8ca1;
        state = 128'h4277_c8b6_b9ca_74b7_d89c_27c2_871a_5ff2;

        #200;
        key = 128'h928b_d84c_5eb2_c366_ae28_f03e_a8b2_aae4;
        state = 128'hab77_cb85_500b_567b_52e7_2374_ad85_6627;

        #200;
        key = 128'hb748_f141_170d_936f_78ee_867c_66ce_627f;
        state = 128'h4100_18d0_0d94_6bca_8ec9_3ff9_4a65_f41e;

        #200;
        key = 128'h1e4d_e54b_471e_24a5_96e3_9350_4321_0625;
        state = 128'h7579_73a9_669e_ec89_e8f4_982b_4435_8ea0;

        #200;
        key = 128'h9462_7e06_c680_c22b_0424_d8ae_8b8b_610f;
        state = 128'h5eab_a8f5_edd7_2450_8998_bcb8_51f4_e9fd;

        #200;
        key = 128'h5c73_9c9c_8111_826f_db20_98de_a865_0a05;
        state = 128'h14b5_56f9_cd16_26f0_c8ba_8811_ed8b_2bdf;

        #200;
        key = 128'haee0_661c_7c75_89e0_1745_84d4_c103_6039;
        state = 128'hdfe4_6c70_cada_a1d5_a047_2823_33a0_5348;

        #200;
        key = 128'h37c5_cc71_172c_c7b3_d497_4a20_1f20_236d;
        state = 128'h02db_71be_b971_3810_38c0_7df1_3a01_63cd;

        #200;
        key = 128'h0b7d_8a62_e65d_40b7_1dc9_a9a0_ed64_07a7;
        state = 128'hb402_476e_1c0a_b118_66ff_1a2d_ebeb_6eb0;

        #200;
        key = 128'h90de_ab3f_37ad_c7fa_13b6_d3df_4423_e650;
        state = 128'h2789_a22d_ced2_0603_6b86_cf97_9282_736f;

        #200;
        key = 128'hc4cb_3f11_4a9c_6a9d_b58f_9437_9862_b64e;
        state = 128'h1188_360b_8f1b_747d_2903_a0e0_80bc_dae9;

        #200;
        key = 128'h0791_794f_ddfd_ed86_f1e4_4065_4d60_fa3a;
        state = 128'hc903_26cc_f4a4_72c4_c482_2e2b_d975_e69b;

        #200;
        key = 128'h81fb_38fa_d045_b2a3_4a06_a9f9_9861_9437;
        state = 128'h1626_c16a_74d4_4280_1ff8_df24_3414_2640;

        #200;
        key = 128'h2529_3392_9f21_be3a_a82e_ed1c_03c4_8010;
        state = 128'h1d0e_f228_2935_d221_2134_5269_3072_a007;

        #200;
        key = 128'h9183_3ef1_1d7f_fc73_ff23_e5ad_f20a_ecb2;
        state = 128'hb67e_2690_78b8_461a_5c9e_b053_2691_74f6;

        #200;
        key = 128'h56d6_fd61_80d3_4886_c669_1aaf_9fb7_ec73;
        state = 128'h180d_97ed_6e0c_e70a_634b_6405_a54f_5b08;

        #200;
        key = 128'h7e2c_b08d_f678_71ea_e61f_9376_290a_d734;
        state = 128'hf2ab_36ab_0c6d_2dfc_fcef_cae0_290f_66de;

        #200;
        key = 128'hf7e7_26ee_6f25_cfbe_cf47_a77c_c39c_2382;
        state = 128'h79d3_8a82_aa8a_212b_aeab_86e3_dde7_860a;

        #200;
        key = 128'h1db6_eb38_ba80_2cd1_5c14_ce9d_9b71_baed;
        state = 128'hb673_b009_b1d6_d5ed_8c08_562b_14b5_dbce;

        #200;
        key = 128'h1bba_8a7a_e495_b61c_2cb0_c352_19ef_53d8;
        state = 128'h8ec8_7516_a83c_efd0_5c11_5278_0b0f_eea6;

        #200;
        key = 128'h471c_f5df_e64d_f0ed_ca26_0bac_8987_67ef;
        state = 128'h00bf_e196_c4ac_ec61_b8ef_1871_5398_bf65;

        #200;
        key = 128'h7614_3f5e_ef35_69b7_979f_4912_638b_3253;
        state = 128'h2f5b_d72a_399d_6028_ebaf_c04a_ada2_06f5;

        #200;
        key = 128'h78ff_d211_72d3_6a43_a2e6_ce04_48f8_0ff2;
        state = 128'h6306_3283_1ee4_07a9_318a_950e_a41e_5430;

        #200;
        key = 128'h88f6_03b0_aeab_4a9e_f6f5_1a41_a561_6abf;
        state = 128'h78c4_dbae_636d_86fa_0cb4_7351_a9c0_d850;

        #200;
        key = 128'hd32a_95b7_c504_979a_3f15_8a5c_ddb7_7a7f;
        state = 128'h44e0_1173_6236_460a_fdd6_201d_3485_e086;

        #200;
        key = 128'h6e18_a454_d3a5_0ad2_c5b1_f25e_7212_84b8;
        state = 128'heaae_c639_3f72_2489_ebd5_e19c_39d0_62c3;

        #200;
        key = 128'h708e_3314_f79e_5b8d_91be_2d3f_beea_37c0;
        state = 128'h3ed0_28e8_b971_6cdd_f5c7_70ea_3006_09bf;

        #200;
        key = 128'hf8c4_9466_5ab2_bfe0_8007_539c_1906_8a3b;
        state = 128'h38c1_e903_bfd4_cdf4_8fb8_a8e8_44b7_eed3;

        #200;
        key = 128'h0356_baf6_f53b_7b8a_7de4_de0a_12c4_6232;
        state = 128'hf3f5_0e8c_2e26_b31b_3124_17a1_4759_f9a4;

        #200;
        key = 128'h4dc3_3d27_55d3_59b9_10ac_b737_a42a_5b86;
        state = 128'h6f50_7329_d054_cb46_0cef_ad8f_34fa_49fd;

        #200;
        key = 128'h57cf_c23b_9d96_a709_6670_4ff5_15b3_ca2b;
        state = 128'hc805_8d5d_0345_d879_d6a2_dea4_2d93_461b;

        #200;
        key = 128'h5c63_56f5_d3e1_9799_653d_d7a6_f7fb_b226;
        state = 128'h19a5_3e95_2f20_49bc_bd74_b0a4_b4e2_417a;

        #200;
        key = 128'h0670_b65f_d069_39c2_876c_9816_5ed8_bc40;
        state = 128'hd945_ad48_ab21_383a_6922_ddae_4f3a_3082;

        #200;
        key = 128'h480f_7904_9706_be46_3c9b_f406_4a8f_a931;
        state = 128'hf01c_7766_0bb1_eccf_6a53_c8f1_83c7_7f3f;

        #200;
        key = 128'h6970_c060_479a_5622_d089_0be7_f8a8_4d02;
        state = 128'h3428_9f87_71a6_25e8_c025_509d_c9ec_ccba;

        #200;
        key = 128'h20d9_50b2_a540_65ba_9e68_f21d_b064_1a74;
        state = 128'hcc06_4aa1_4d22_4db1_522d_34a5_6e16_d0f2;

        #200;
        key = 128'h4f1d_8a4c_cbd5_b8a0_298b_50a2_3484_b97b;
        state = 128'he085_2ccd_9d47_ba42_db1b_f8fb_6799_e26a;

        #200;
        key = 128'h17b6_e1e8_a70d_6cb2_bc72_2fe4_923a_991b;
        state = 128'hd956_a21c_35f3_506b_1b9d_9364_2211_59ad;

        #200;
        key = 128'haccc_2048_f01f_9d4d_c538_ae0a_2f26_e57c;
        state = 128'h93ae_2181_d708_3efa_4ea8_8dca_af85_1e8b;

        #200;
        key = 128'h420f_4acd_2ec2_71d1_ef71_ec89_8d71_1b8c;
        state = 128'hcce2_efc2_31a8_f829_8249_0aa2_117a_fd11;

        #200;
        key = 128'hcde3_5585_f938_7ca9_e5d5_fc61_04a5_1bd3;
        state = 128'h4f33_502b_5ac7_76ff_4070_20da_20af_ed8b;

        #200;
        key = 128'h1373_bc00_5c1c_9b50_ae15_08ea_3851_534b;
        state = 128'h76a7_b650_1058_5692_c96f_87dc_f92d_580f;

        #200;
        key = 128'h0185_cb54_4412_f831_2c82_d952_e28a_ca83;
        state = 128'h68e8_1950_9eb9_1e7a_884b_d355_730e_beb7;

        #200;
        key = 128'hf6f2_5e50_03ff_72a4_688c_1db0_30cf_1d7f;
        state = 128'h2a38_a4e7_b90e_119c_583f_337d_e420_f367;

        #200;
        key = 128'h5a9f_45f4_0f35_efb9_d03b_4beb_73bb_4b17;
        state = 128'h8d85_70cb_ff8a_faad_a2a4_75c4_0647_af66;

        #200;
        key = 128'h6857_55ab_207f_440f_648d_c20f_9fdb_b1bf;
        state = 128'h264b_fce9_f29a_f3dd_c4e5_746e_47ee_a3f6;

        #200;
        key = 128'h4a47_4f81_44f0_271c_983a_761e_fa8e_7edf;
        state = 128'he6e4_9560_969b_c2c2_21dd_2776_ba8e_14d4;

        #200;
        key = 128'h53b7_fce7_fe40_533a_9bdf_f0d9_4d30_59cf;
        state = 128'h3d2d_908f_2b7f_7508_f2a1_e684_3c3e_1a6d;

        #200;
        key = 128'h138a_0a2b_9105_cbfc_a05e_1e57_f926_81b2;
        state = 128'h5db1_6e40_ea5d_6519_6eb9_e64d_f5fa_d682;

        #200;
        key = 128'hc1a0_18b1_123e_aad1_935a_9da4_8c22_a03a;
        state = 128'h3c51_f43e_6a9e_718d_d43d_4751_51ce_058e;

        #200;
        key = 128'hd436_ea52_27a0_0f58_6a73_9814_7da7_bf82;
        state = 128'h4de7_a3fa_1778_f20d_1c8e_b5cf_5093_8e14;

        #200;
        key = 128'h53dc_76a2_4007_12a4_32c9_1bb5_86f1_653a;
        state = 128'h584e_a524_aae4_4a6f_a618_2ba3_7d6d_e1c9;

        #200;
        key = 128'he86a_2a30_b9c4_bebb_0105_8b76_05a9_0888;
        state = 128'h24e7_26af_f0b9_ebd4_ce32_733b_7632_50cb;

        #200;
        key = 128'hba87_3a54_c491_d1de_f3d8_2a7d_d311_3bf5;
        state = 128'h0383_3383_2ac2_5fd3_941d_63d8_477e_3b3c;

        #200;
        key = 128'h472c_1729_8e24_063f_d27b_77a1_95a5_586a;
        state = 128'hb7d3_2167_3c6b_dca9_2445_6c5d_eeae_8366;

        #200;
        key = 128'h70e9_cbaa_8f1b_fb3f_6009_44a0_9b42_24a4;
        state = 128'h3f6f_4b36_2f86_8fda_4df8_a5af_41a9_598a;

        #200;
        key = 128'he128_2b98_2834_5c79_a9b1_1b6a_0bd4_3355;
        state = 128'hef9e_2d08_429c_0f3f_1b52_a96f_f1e2_70b7;

        #200;
        key = 128'h4062_bef8_6090_f566_7b1d_907c_99a3_9e5e;
        state = 128'hae4e_2a4b_d048_980c_7bc8_03c3_08eb_00b4;

        #200;
        key = 128'hc636_1082_b89b_2305_7bfa_0489_7bf0_4aca;
        state = 128'hb92b_63e4_8f18_5612_7ee1_da20_8fa3_662d;

        #200;
        key = 128'h2841_c25c_e555_8c22_d176_fb5b_6ad8_e607;
        state = 128'h6cb8_7943_2d12_35ea_2eed_a5fe_56a3_629c;

        #200;
        key = 128'hfeb6_bf6e_a648_e144_c059_d266_e820_6d62;
        state = 128'h2de9_d829_0c3f_2f69_7260_7d2a_85e1_451d;

        #200;
        key = 128'h56ab_0e18_1615_555c_a3c5_6f75_c642_1cc3;
        state = 128'he5d0_295f_6b61_4919_e0f1_af05_bb27_4d11;

        #200;
        key = 128'hfbc8_c2ee_e67f_d563_6c75_1fa2_9d7d_877b;
        state = 128'h180a_df9b_dbd2_7131_8cbb_4c3e_954e_3361;

        #200;
        key = 128'h098a_cd81_448f_1cf6_a14a_b09c_3c84_83da;
        state = 128'ha21c_85a8_2e34_0ff7_074e_53cc_90cc_bc69;

        #200;
        key = 128'h4ecc_265c_75d8_5934_c97e_7d8b_c947_1c86;
        state = 128'hec89_2e32_737a_1264_d445_8256_b60a_4cc4;

        #200;
        key = 128'h38a4_66ce_adf4_139f_217c_7eb9_dad6_9c6a;
        state = 128'hb933_f43a_bf01_02e2_a90b_8e2f_f858_9c50;

        #200;
        key = 128'h2341_94cd_0412_0c37_27f8_1185_25ac_be78;
        state = 128'h5d89_19a1_544f_1169_d1de_ae4f_db34_51f1;

        #200;
        key = 128'h165a_9a4c_9aae_ef89_2ea2_d40f_482c_66eb;
        state = 128'h43f6_ce00_8f14_6936_51dd_18e5_10ea_ce06;

        #200;
        key = 128'hf994_c798_b6a2_acf9_c54a_2d30_7d96_deb6;
        state = 128'hd6f2_6d30_39b7_aa33_d40a_e2d7_63aa_d74f;

        #200;
        key = 128'h32cb_bddf_7b34_2172_b8de_f027_0373_8b23;
        state = 128'h33af_5521_9867_3c6b_e171_af39_9c81_d6c1;

        #200;
        key = 128'h0b9c_f6d0_71ca_007f_5a92_f0b1_b501_12f8;
        state = 128'h1177_a323_c7a8_3b8d_283c_bf54_1537_a0db;

        #200;
        key = 128'hfbff_0683_b776_89fa_07f4_e1d3_51a8_b477;
        state = 128'ha439_e2fe_f86e_0413_ff9c_61f8_8626_e17d;

        #200;
        key = 128'h12a4_3f31_76db_4108_d9df_f5d8_bf4e_dc1d;
        state = 128'h0228_c4cd_c87b_ed0f_55ea_8048_9a8b_a33d;

        #200;
        key = 128'h58ae_df77_0161_19ab_3ae5_2ee8_71b7_a517;
        state = 128'h0c61_4466_0538_d4d3_1124_3bdc_f9ee_35df;

        #200;
        key = 128'h6e01_6c25_143c_7d59_1ddb_d344_69e7_94f9;
        state = 128'h7a83_f488_c692_4ddc_37b1_c43f_cd61_425c;

        #200;
        key = 128'h634f_3e40_41f5_f59c_6f5f_b1e9_bda1_bbcd;
        state = 128'ha917_915f_4f4e_2534_e1a0_b180_0cbe_bbaf;

        #200;
        key = 128'hceeb_b70b_544c_8ae4_dd4f_e239_6477_2a26;
        state = 128'h29d0_0e94_fe53_dc93_ce25_fe20_e29f_59f3;

        #200;
        key = 128'h5886_370f_3d8a_8904_53da_8ac7_6242_396e;
        state = 128'h0f02_8cae_51f0_a12a_593b_7847_0731_8941;

        #200;
        key = 128'h1918_5d16_4236_db2d_d6a4_2d0a_eb8a_659e;
        state = 128'h6b99_6487_9c55_c007_7283_251d_56ae_d8f5;

        #200;
        key = 128'h1664_bc0f_5fe9_c875_5e92_149e_6af9_2070;
        state = 128'h63da_6dae_5946_6030_56bc_27c1_1fa9_c684;

        #200;
        key = 128'h23bd_b17a_9e1a_e5de_da08_7d2e_2414_16fd;
        state = 128'h02d7_b80a_ba69_5b7a_845a_2d81_bc1a_bf2b;

        #200;
        key = 128'h33af_1ef9_cd6a_2d53_d94c_2b60_08cb_4da2;
        state = 128'heaae_ebb1_4334_0a11_d0bb_f28c_ce15_7fe8;

        #200;
        key = 128'h0ed7_2e12_24e5_e0cb_4e57_ee1c_828d_8085;
        state = 128'h5def_4711_7b57_ea2b_58a8_1a4c_5b10_af5c;

        #200;
        key = 128'hb91e_854b_7027_88ff_1622_b3c7_6d8e_dabe;
        state = 128'h7c15_10bc_bbf7_7f56_dfa4_4fdb_c760_7aa9;

        #200;
        key = 128'h3c6e_0c3e_6180_a42a_3f7a_6ff3_cfa1_c7d6;
        state = 128'hf590_c152_d5ff_0756_886b_d1e6_a590_d121;

        #200;
        key = 128'ha77a_a27c_0632_91a3_a43a_fbfc_948a_7d6c;
        state = 128'h24e3_035b_d1c9_5dec_dbbb_df3c_d9c7_3ee6;

        #200;
        key = 128'h1143_090d_62a0_7f12_5058_9b79_dd20_ff43;
        state = 128'h52fb_5583_006a_fee6_5408_0a70_c24a_2891;

        #200;
        key = 128'hb81c_5490_3197_598a_8deb_fe1a_9ef3_19e1;
        state = 128'h02bd_84c2_ec0d_f95b_9967_33cc_aa6d_c648;

        #200;
        key = 128'h0c18_e83a_117d_642f_c58b_8805_8c94_ba14;
        state = 128'hf52e_1aef_604b_9baa_962c_2cce_3bd1_0fa2;

        #200;
        key = 128'h5f15_1068_1ae5_488e_dfd7_6292_1edb_a454;
        state = 128'h30b1_187a_bd84_3a9f_60a9_c663_7399_f53c;

        #200;
        key = 128'hc419_ae17_400f_e82a_c35e_b078_7294_4668;
        state = 128'he924_7d03_5d50_1c01_cffd_bc58_a325_dce7;

        #200;
        key = 128'h8224_d1ef_1b2a_dc14_ee83_dab9_aa3b_fea5;
        state = 128'h9d9c_abcc_4fbd_d3d5_9a4f_db84_6d5f_7336;

        #200;
        key = 128'h7550_162b_3f4e_3129_aa12_53ff_d742_998a;
        state = 128'hc15c_c020_c1cc_0861_9fa3_0035_1781_3ede;

        #200;
        key = 128'hd139_0943_913f_a3d3_2276_246a_a592_b35f;
        state = 128'heaf0_b068_3e11_5d43_ac55_d099_c972_79d2;

        #200;
        key = 128'hbdf3_26ce_d7e2_62d4_bcb1_4cfb_a1b5_f059;
        state = 128'h033a_6493_d7b7_834b_fe50_4f87_54d1_fd46;

        #200;
        key = 128'h3101_9897_f680_afd1_731d_07a0_4765_1544;
        state = 128'hee28_f02d_a18d_c222_131c_b516_df92_7683;

        #200;
        key = 128'h895e_4b15_a62d_39ae_25dc_55c2_89ad_e5dc;
        state = 128'hf0cd_034a_3511_da1c_9f5f_1019_763d_c8a0;

        #200;
        key = 128'ha8a3_685d_2687_cecc_2e07_f137_471c_4cb9;
        state = 128'h82cf_0f0d_b475_6602_b3b8_5026_7877_d48d;

        #200;
        key = 128'h1bb4_67ba_cff1_99ba_b16d_34d1_a2a1_4b92;
        state = 128'h8004_01af_eec5_7e50_c524_9c33_9769_6509;

        #200;
        key = 128'h285c_86a4_fb33_dec1_f684_af86_30eb_568a;
        state = 128'h122c_1252_2e63_d309_51a7_0025_8638_030a;

        #200;
        key = 128'h1902_8a81_a2e8_30e1_b923_0a02_672b_f2fd;
        state = 128'hf74d_2be2_5867_c052_e937_5720_c527_95be;

        #200;
        key = 128'hee65_2f52_88a1_6ac4_9bd1_8dff_e771_2c02;
        state = 128'h511d_8d02_4371_dfde_fa0a_f301_bdfd_d0bc;

        #200;
        key = 128'h98b6_2381_1e5f_8c44_185c_a814_620e_bb0e;
        state = 128'hc5aa_b28a_4e98_ff06_a835_4c36_8dc7_1fcc;

        #200;
        key = 128'hf3c1_022b_3f05_dbda_5829_6d0a_dbef_2e8f;
        state = 128'h5980_3e3b_19a5_65eb_8dda_a15f_a88b_0e7a;

        #200;
        key = 128'h80d6_d8f2_90e1_8406_7ec7_81ac_7171_3704;
        state = 128'ha7d1_38a3_1d69_96d4_9855_d35a_38c2_78d2;

        #200;
        key = 128'h4b5b_db1a_c39b_1d83_5e3c_242a_abf7_905a;
        state = 128'h1ca1_27ce_89a5_7dd8_65fd_80f4_6dbb_a9d7;

        #200;
        key = 128'h0c8a_15f0_0498_135b_c023_ac79_43f1_edd2;
        state = 128'h384c_14f0_8781_ea5f_7033_e5b3_c19c_9728;

        #200;
        key = 128'h99e5_d57a_efee_778c_cbe5_2e38_a302_9cf6;
        state = 128'h54fa_766e_a254_4be2_7325_66b3_c828_619b;

        #200;
        key = 128'h8cca_cbc5_8518_bd88_2d32_b765_40ff_27e6;
        state = 128'h535e_0952_6041_1581_89a1_5fc6_5799_4de5;

        #200;
        key = 128'hd832_ade8_0fde_5f0c_fc9f_ecf4_e472_05d9;
        state = 128'h5f30_ce6a_3031_a74a_e7c2_b549_891d_112c;

        #200;
        key = 128'hbe53_702a_7820_574a_4439_eaa3_04b2_9e8f;
        state = 128'h5a1d_ef56_45a5_7374_07aa_46e9_9fbb_7c2f;

        #200;
        key = 128'h749c_59fc_c22d_601d_34fa_11c3_7c32_5c0c;
        state = 128'he5f2_c147_38ae_ad4e_ef8d_be03_7743_ab84;

        #200;
        key = 128'hbc80_8662_f452_940d_3cf2_a075_6098_002d;
        state = 128'hd266_c5e3_2c0c_451c_93fe_c1ff_2b67_0be3;

        #200;
        key = 128'hbdbd_88eb_3765_5f91_6fd8_21ec_4929_aa18;
        state = 128'hfe8a_9904_d40d_65bf_8fe9_384a_cb97_5f59;

        #200;
        key = 128'ha5c6_ea95_99b6_887f_cb04_9075_9d15_99c9;
        state = 128'h74d4_fb41_8efe_1d01_ce35_48b5_62ba_b118;

        #200;
        key = 128'h21ca_714a_1a4a_8865_5274_477b_067c_f12b;
        state = 128'h7049_28c4_aff3_31b7_9378_c6ce_69c4_1561;

        #200;
        key = 128'hb6cf_1b5c_71e4_e1bd_8410_55b6_18a4_320b;
        state = 128'h3a51_fa46_0d84_b7f9_1326_fef1_c4f5_cf5e;

        #200;
        key = 128'h4866_b4b7_2431_841e_1b77_1e30_eab1_7f5b;
        state = 128'h57e7_618b_6772_499d_8ce4_2c8e_7113_0f6c;

        #200;
        key = 128'h4e98_6616_f573_68a0_e13e_e654_3289_1205;
        state = 128'h07ba_2372_6bd8_fccc_05f9_fdd8_1d2b_1fd4;

        #200;
        key = 128'hb226_9b43_0247_868c_5809_8509_0f4e_6c6d;
        state = 128'hfbaf_0c9d_27ec_7ce8_daf5_6dd1_a260_a0f3;

        #200;
        key = 128'h7981_29cc_ea34_af41_ae9a_122e_69a0_2340;
        state = 128'hab8c_0d85_c11d_e32e_6117_a881_d56e_e7ae;

        #200;
        key = 128'h58c2_1def_28fe_8ac3_13ae_1d15_b4b4_d20f;
        state = 128'hb02e_879b_05df_1af3_0557_31bb_df78_b119;

        #200;
        key = 128'h5b52_b865_c873_1230_211d_c1e0_0b53_bae7;
        state = 128'he418_07ba_2a85_8cb2_49a3_b606_3019_c5ae;

        #200;
        key = 128'h0bff_7f30_729d_652f_f9bc_7c9c_d2a2_1af0;
        state = 128'hb7ea_a790_ed6d_aeeb_b2a7_c9c0_1674_ac55;

        #200;
        key = 128'h923a_18a0_165f_16cf_a0d1_6810_e229_69f0;
        state = 128'h7e95_210d_78dd_a363_29dc_edb5_2ca4_9e35;

        #200;
        key = 128'h7289_b85e_5e80_b33d_4d62_3e58_8e94_1f3a;
        state = 128'h3405_276f_cd8e_e65c_9c20_f197_9702_17e7;

        #200;
        key = 128'hb35e_df4e_1cf6_8b85_e3f8_2c3a_62b5_c801;
        state = 128'h29e7_242b_b464_59d6_c9ef_5496_ae66_68be;

        #200;
        key = 128'h9391_b219_b723_1d0a_d878_0983_5311_bf44;
        state = 128'he9af_40c8_a2d5_9ee6_30d8_4827_97e3_968f;

        #200;
        key = 128'hb79a_f807_6293_2b75_c9bb_ed86_4c66_d489;
        state = 128'h84f7_ee79_f3fa_bba5_c6e9_9eac_c14d_ee37;

        #200;
        key = 128'h9b79_5631_bcb5_03a9_1d3e_3630_e23c_b634;
        state = 128'hc788_9bc0_85cd_bdab_7fa8_39f3_4de0_d674;

        #200;
        key = 128'h1eb0_cadd_55c9_8a8c_53a5_a266_d1d1_e005;
        state = 128'h75da_1a33_39ce_161a_51d9_3a4d_2cde_6b66;

        #200;
        key = 128'h7015_a571_4160_4106_f24d_67aa_2183_25a8;
        state = 128'hf715_4cc5_6a6b_b652_9ac3_3ea4_87db_4be0;

        #200;
        key = 128'hb55e_919a_ed55_460f_f3ac_2817_097f_bd3e;
        state = 128'hea45_09f8_acc2_7a88_eb68_3f0a_2b16_d61d;

        #200;
        key = 128'h7623_0c38_c9ab_4e62_5a2b_4d1e_b691_9075;
        state = 128'he4d4_cbed_0938_bd50_44a2_43d5_96ec_a2da;

        #200;
        key = 128'hb7c1_c9a6_5ac1_96ab_5753_38ba_b13e_5ca9;
        state = 128'h3c0c_1d75_61e6_85a7_cf25_7b35_e071_03b8;

        #200;
        key = 128'h8c3f_423a_0067_41e3_14b7_e7b9_9a3d_aed7;
        state = 128'h496b_a183_76b1_a552_448b_629f_f678_b87b;

        #200;
        key = 128'h36a9_a369_c69f_871d_c6b4_b5a6_00a1_2041;
        state = 128'hd6d6_16c0_7ba0_ad6e_b020_ea83_ca00_2c43;

        #200;
        key = 128'hb9bf_afaa_6634_7188_b0fb_d407_f245_f61c;
        state = 128'h18b0_04b0_30a3_fa7d_d7b2_5b34_f711_1b69;

        #200;
        key = 128'h9012_15af_534f_3b3f_3c35_5a5e_cbc9_8e51;
        state = 128'h27fe_39c6_450b_2b71_07d0_76e8_5c16_2a2e;

        #200;
        key = 128'h8fa6_824b_7965_6491_4b65_ef92_0085_b9ce;
        state = 128'haaa1_a4f4_ae49_6a79_33fa_18eb_98bb_b8ed;

        #200;
        key = 128'hb972_a922_41b9_dd46_c94d_0d36_d2f9_a5c8;
        state = 128'hd085_219c_7ca4_d409_7af7_2069_3556_4cfb;

        #200;
        key = 128'h744c_f14c_26c2_669c_c5a3_fc41_3f6f_b097;
        state = 128'h51a5_2b90_5d26_f7cb_e3bc_5478_7c67_0871;

        #200;
        key = 128'ha3d3_50be_8650_1e3e_a226_10f8_4cdd_2159;
        state = 128'hd391_8d51_d81b_235f_cb14_1fe6_0036_36c5;

        #200;
        key = 128'h1023_22d9_2916_22fc_261d_9653_6796_c6b0;
        state = 128'h053e_6b26_e21d_1ea5_3eea_1877_2cda_2fc7;

        #200;
        key = 128'h11b4_7a11_b8bf_ebe6_c54c_587c_9fb0_b6ab;
        state = 128'hcffc_ecff_c994_fe58_d04f_c86c_8c42_04bc;

        #200;
        key = 128'h7b1f_9719_2b48_9a8c_ed8b_a320_7894_d683;
        state = 128'hd0ac_4aaa_a803_8590_0aff_8e66_8958_2d49;

        #200;
        key = 128'h4915_0995_4204_ace5_3fe1_af10_2117_b4e9;
        state = 128'hd417_68ff_4c38_16f4_4c77_276f_6242_1559;

        #200;
        key = 128'h408e_f15c_8bed_99b4_4cf2_ca0e_bfc6_6ff7;
        state = 128'h7190_0595_5846_39cb_2486_e794_90c6_8cb4;

        #200;
        key = 128'h317b_a584_2e9c_01eb_1f3c_b3b4_22cf_fc6e;
        state = 128'h386b_3f98_4811_dfb4_2d5c_f17f_218b_094b;

        #200;
        key = 128'h36ab_3f9d_2a4f_d613_9872_bafd_d16c_d08b;
        state = 128'h15a8_c0ec_7e94_cc98_a50b_b96f_2d70_779f;

        #200;
        key = 128'h1fbe_043f_f60f_f4be_3ff0_50d2_e424_3189;
        state = 128'h966c_581f_030a_dd8b_8a13_d4b7_43c7_a62f;

        #200;
        key = 128'h6e8c_9941_7a7f_45bb_97b4_49b9_9455_4b0f;
        state = 128'hda6d_1466_4d07_1589_32c9_195b_5c02_7d18;

        #200;
        key = 128'hfd44_2a90_6330_4640_271c_d5f7_3e6d_8439;
        state = 128'h2806_09fd_74ea_c565_3a54_01bc_cb68_7416;

        #200;
        key = 128'h6d59_5c81_95d6_3780_c769_0b1c_fde2_f2cd;
        state = 128'h1a27_3c39_95ff_9192_7538_1133_982d_b9e3;

        #200;
        key = 128'hcbfa_7ebc_b5ef_2100_db92_865d_3367_b037;
        state = 128'h4dd4_869d_5cee_0339_1d2f_e57e_64d9_941a;

        #200;
        key = 128'h58ab_a885_9f76_5a49_6b43_79a5_cb88_fd84;
        state = 128'h9a3d_939e_a00a_3fe7_22b6_8f8e_c0eb_952f;

        #200;
        key = 128'h2bea_21ff_4be0_4945_732c_3653_e609_f31f;
        state = 128'h62a9_7753_37ea_3f60_27db_1533_3267_553d;

        #200;
        key = 128'h7d6e_4f8c_440e_b339_659b_95c9_d5ce_7007;
        state = 128'h19d5_748f_15f9_7b42_7d74_6eda_ec01_b3f2;

        #200;
        key = 128'h3e9a_8e8f_d904_460c_c1e8_e7c7_2a6f_dbfb;
        state = 128'h0678_da0b_06fb_d2c8_c159_121e_fef5_2a09;

        #200;
        key = 128'h0b91_8521_b460_c5f0_f4e8_3085_d2f6_6118;
        state = 128'h4ac0_b0c9_73b3_8281_8636_90ba_02f8_7c17;

        #200;
        key = 128'hed5e_aa0b_cd70_1fd2_dbc1_3a74_5dc6_6f09;
        state = 128'hee8f_88ea_d3c5_ff87_05ae_50ab_16f6_7616;

        #200;
        key = 128'h58ca_2921_af82_0bd7_0f4a_a60d_f133_7dcf;
        state = 128'hc0e9_44b3_a39c_14c2_baac_f27b_7f08_3e0c;

        #200;
        key = 128'hf3c4_6f2f_dc89_e55f_88b7_594e_39a7_9317;
        state = 128'hbb5b_51ec_2fc3_2150_6187_2bd0_7dc8_89a7;

        #200;
        key = 128'h3b61_bab2_e0d8_47f9_dca1_e0bb_68ba_a907;
        state = 128'hd20f_c360_34c9_769b_8962_96a3_a18b_0b0f;

        #200;
        key = 128'h0ef2_a46d_4b13_8579_fc2e_6e3f_abde_faae;
        state = 128'h8e82_aa05_4cc2_2b60_bdca_7582_ef12_eb47;

        #200;
        key = 128'h4bbe_ee50_fb1f_861f_f36e_072f_5dd3_9783;
        state = 128'h5e60_76f5_3c83_dd6c_2a83_8b7b_bc83_125b;

        #200;
        key = 128'h30c4_f497_9bfd_f1dc_8933_55d9_c424_5cf3;
        state = 128'h0bdf_e479_b4fa_aed0_8c98_d64e_017f_bb8e;

        #200;
        key = 128'h5d14_e0c5_722d_4b2b_907e_9aca_67b6_c7d8;
        state = 128'h2ab1_a09a_0e50_e476_ee4b_0424_8dbe_98b6;

        #200;
        key = 128'he6c8_c7a7_1151_2ee5_d297_0fa6_4cdb_ff1a;
        state = 128'h9abb_b020_87b5_bfd7_1aa2_62a2_c4b8_ed38;

        #200;
        key = 128'h8c4c_3d75_33b7_febe_5f4f_bea8_6f52_dacb;
        state = 128'hd8d3_8632_4d81_ad10_5376_afbe_a469_a72a;

        #200;
        key = 128'hbf03_827c_4718_48d4_ca44_bbfd_a60a_62c6;
        state = 128'h73df_4914_531a_7410_d883_ff05_77b2_d0db;

        #200;
        key = 128'h5c8a_7728_d511_d595_f628_7ec3_9641_5f8d;
        state = 128'hdffa_949f_6f10_53f3_03c9_9bec_01b0_4817;

        #200;
        key = 128'hd9fd_0960_d04c_4986_0646_6ff8_7b20_6cb6;
        state = 128'hf07d_ac55_dfde_c16e_6a5c_a82c_de40_ad34;

        #200;
        key = 128'h2ab3_14e0_f104_51f2_9149_649e_353f_2625;
        state = 128'h5c32_0c75_7689_94de_54bc_35e7_95d2_501f;

        #200;
        key = 128'hc7a5_fe0e_8680_51ff_77fe_d0a7_6672_97c1;
        state = 128'he7f3_41f3_1880_fa0b_cb69_e07b_f397_0f4a;

        #200;
        key = 128'h8d2b_86a9_4227_e01a_67f0_8cfb_8c30_d053;
        state = 128'hfd0a_d94a_bf78_9266_6ea4_2d05_cda7_752c;

        #200;
        key = 128'hd2bd_6235_8b09_acc7_0f7c_ef62_b0da_5379;
        state = 128'h5f3e_b9e8_b28c_99f5_c1d1_23e7_28ad_7878;

        #200;
        key = 128'h4429_4071_8be2_8905_9f17_10f2_3f85_98d5;
        state = 128'h3045_6b62_62e9_5428_b92c_41ba_faae_d32d;

        #200;
        key = 128'h9e97_3322_2261_7854_40c7_74c1_d54f_3978;
        state = 128'hd4e4_0415_e0e3_9a3b_caea_82e5_1aa9_35e1;

        #200;
        key = 128'h31a7_84e4_c7b5_1608_b199_23f9_0b08_216f;
        state = 128'h3b96_7d05_e9a5_da21_34dc_3cba_828e_39f6;

        #200;
        key = 128'h3e03_dab3_983d_3c0f_f3d4_e361_63b5_3539;
        state = 128'hd6c0_67e6_1307_a0f5_2254_a136_de70_544a;

        #200;
        key = 128'h3b50_cc52_0ced_8964_c77e_f07a_e883_8836;
        state = 128'h49a7_64be_02cd_4d11_63d9_d254_d3ba_8524;

        #200;
        key = 128'h9dca_2836_164e_c64e_950a_c174_bd9b_0813;
        state = 128'hbb1b_133f_633f_0f79_f0ed_06f4_8627_b914;

        #200;
        key = 128'hdc4d_3ad1_7a8c_4ad8_22d3_ab86_f091_286c;
        state = 128'h5a97_1bb9_fee7_758f_34b0_1eeb_6e9f_390d;

        #200;
        key = 128'hf122_a380_3411_e976_a917_bfd5_3263_2e76;
        state = 128'hc221_5879_4e32_f0b3_40be_967b_a19c_eff8;

        #200;
        key = 128'h3072_ec95_7d2e_97bf_9243_b685_4385_ddfb;
        state = 128'h904c_6a8a_9241_4484_1478_670e_7240_e87f;

        #200;
        key = 128'h46eb_ba7f_51aa_83f8_8dbb_168d_73ce_676f;
        state = 128'h3b16_2adc_6369_2857_6ffe_b794_9218_d90d;

        #200;
        key = 128'h6519_e012_30b4_6f35_f7b4_b5de_bc24_c1ad;
        state = 128'h826b_6da6_5b04_9a4b_4f87_1977_ffd3_6940;

        #200;
        key = 128'hc33f_5f54_454f_0a10_73bb_f102_976b_e788;
        state = 128'h960d_d6e3_427e_c3d6_0749_b256_7bc1_dbf3;

        #200;
        key = 128'hf214_dc82_7143_f0cb_a4c4_2197_746f_3c2a;
        state = 128'h2644_bb2f_f983_63cd_1315_18b9_2ae8_d8f8;

        #200;
        key = 128'h2224_6641_1b8d_7be3_62f3_6cb0_07b5_bcc3;
        state = 128'h73b5_d1be_46a6_f96c_4dd7_4c45_d737_c18c;

        #200;
        key = 128'hd433_138d_ade4_f592_57a2_eb81_5a8f_1b7a;
        state = 128'h44cd_4185_3883_aa0c_7d14_de48_cad0_6f9d;

        #200;
        key = 128'h68a1_ef0c_cb2b_ca9b_2dad_f3e0_4813_7df3;
        state = 128'h5d83_370e_4e5e_565f_8e21_1d1f_bc32_3dca;

        #200;
        key = 128'h211a_75c9_cde3_e96e_26f2_edb1_fd8c_3889;
        state = 128'he926_8d99_71b7_1443_1ddc_e328_d032_1c1b;

        #200;
        key = 128'hd5fa_c0f9_2027_76be_72b0_169b_7524_1ecd;
        state = 128'hc3cd_8322_ec72_bd88_34df_8fa0_c89f_638f;

        #200;
        key = 128'h4403_a79e_fd6a_07ba_40dd_17d9_013f_6f47;
        state = 128'h9ead_a30a_6645_350c_b07c_6dbc_3ed3_9f77;

        #200;
        key = 128'he9e7_2f13_7339_d163_162a_4cef_0a6b_0b25;
        state = 128'hbcbc_0041_0e9a_d038_c0a4_393d_8e7e_a643;

        #200;
        key = 128'h7b30_a652_9b48_d4e1_2da7_3b9e_0466_e229;
        state = 128'he542_6e2e_fa36_08af_db8f_a358_a81d_b506;

        #200;
        key = 128'hb06e_f04a_74ce_aff0_0a18_ae3a_7823_eaec;
        state = 128'h6fe7_efb0_f8d6_a1a0_7ab0_e17b_51da_7960;

        #200;
        key = 128'hfd44_7f39_8964_de71_241e_5ede_ddff_9c8a;
        state = 128'h545f_2fcb_3402_4540_11e6_1392_7f14_8779;

        #200;
        key = 128'h08dd_71e5_fe6e_4f72_8d3c_3603_6f5a_0300;
        state = 128'he824_257f_0afa_dd37_9137_821f_244e_940f;

        #200;
        key = 128'h701f_4be4_81ad_07f7_273c_44d3_c036_117b;
        state = 128'h5bf0_92d8_8921_1a6a_8fee_88cb_7966_17db;

        #200;
        key = 128'he467_40d9_9ba9_75fd_a6e6_e239_334b_e688;
        state = 128'hb30a_8b5e_871b_f79d_a2e2_ba41_a159_29ad;

        #200;
        key = 128'he04f_b22b_99a8_ae25_fbc9_de6a_0e75_5952;
        state = 128'h4337_8702_e8df_a0a8_d584_2b91_d90d_ea4a;

        #200;
        key = 128'hf6d6_98f7_c039_3ce6_54e0_cbae_035d_a7c4;
        state = 128'hea10_fd2c_8531_1ca9_1983_a098_6903_07d0;

        #200;
        key = 128'h1ea7_50cc_e9c5_4c41_c426_9222_7a93_114e;
        state = 128'h10ca_bc32_38f6_788b_78d1_20a8_24da_61f2;

        #200;
        key = 128'hb88b_9f02_b1d1_fd33_12c2_6379_9333_9e0d;
        state = 128'heed5_eb36_a281_9b34_f20e_8c70_f57d_993f;

        #200;
        key = 128'hb03a_c51c_ba02_dc41_51b0_791c_84d3_1186;
        state = 128'hbba8_7a4d_96b0_1720_f482_e28d_c6de_dc45;

        #200;
        key = 128'h5bfa_d3db_9d64_34f9_a241_ca5c_1665_7c86;
        state = 128'hc931_da36_fca7_18df_3503_1b63_daac_8b8f;

        #200;
        key = 128'h662a_b5f1_8341_6d8a_812b_710a_347c_d112;
        state = 128'h1091_8e37_7440_8757_96e6_3060_0d42_1422;

        #200;
        key = 128'h5008_c4a4_0a18_9ebd_c4ba_3fc9_b5f2_50dc;
        state = 128'he3a6_88cb_08d3_a05d_5083_883a_6f4b_2754;

        #200;
        key = 128'h463a_e4c4_e916_dd1f_813d_af37_6b42_f174;
        state = 128'h5122_b24e_43e7_fe63_991c_b66c_4621_866a;

        #200;
        key = 128'hc770_b5cd_90c6_f5d6_840c_8a3e_42c2_2f39;
        state = 128'h4117_5e3a_ff3c_590f_2166_e246_75fd_78bd;

        #200;
        key = 128'he274_947e_7e1b_3647_5875_ca51_90c9_e8b9;
        state = 128'h9868_1bfa_36ab_b70f_2c8c_4a79_958f_c715;

        #200;
        key = 128'h0bba_bf23_fb98_96cb_1a2b_d7f4_9268_1288;
        state = 128'h7425_1d49_ee7e_d5ec_7376_d47a_5530_2649;

        #200;
        key = 128'h39de_758a_1df8_18eb_2792_6507_127b_faa0;
        state = 128'h328a_bd77_518d_04a6_9d1c_167d_0a41_e33d;

        #200;
        key = 128'h760f_7746_f526_7859_abc0_6dca_2384_d577;
        state = 128'h1dce_2192_77bc_b8fe_d63b_33d1_2453_7b5c;

        #200;
        key = 128'h9f45_7f58_32f1_68bf_8bad_f5db_cbb4_7fb2;
        state = 128'h63b1_456a_a1fe_5bf8_70e9_d916_0e78_a4ae;

        #200;
        key = 128'hbf5d_93b3_d80c_1eaf_497a_3ad7_934c_e464;
        state = 128'hf022_f82b_127d_8af2_0a85_aa96_edfa_71ce;

        #200;
        key = 128'h9729_a208_1359_1fb8_0412_c579_07bd_918b;
        state = 128'hf816_91b9_99c5_1136_39df_f1fc_d7d9_411b;

        #200;
        key = 128'h4c67_a19a_ca5e_1f15_f488_9b5a_5060_3ee7;
        state = 128'hc320_0817_c1c5_5718_de2c_4f6c_cb9b_dfe8;

        #200;
        key = 128'hbef0_4ff2_a135_5f05_6ad7_465e_7563_8f2e;
        state = 128'h363c_d26e_03c5_0e8d_3f9d_0137_8775_2ff6;

        #200;
        key = 128'h5b2c_b49d_e208_84bc_893d_6aca_5ba7_903d;
        state = 128'ha03b_2569_5c54_d794_b719_9690_cf7e_cc36;

        #200;
        key = 128'hf791_9943_5aef_1d5b_396d_ec2c_f067_ed69;
        state = 128'hd20a_8b8e_81be_337e_ac42_6f20_d9fb_098f;

        #200;
        key = 128'h59a3_773d_524d_5b45_a5da_33bb_dc32_82be;
        state = 128'hb791_c622_03cb_67f8_c27a_eede_09e3_08ed;

        #200;
        key = 128'he445_e772_bdba_39cb_7cb9_64ed_96b1_74cb;
        state = 128'h3b57_b6e1_7f97_e6be_d0d4_5414_c1e4_d187;

        #200;
        key = 128'h113c_4eb0_7274_edf1_4bc4_a891_fec2_b991;
        state = 128'h14d5_8797_db32_f7ce_9c4c_ecbd_dae1_38f7;

        #200;
        key = 128'h243f_e0fd_23d3_e22f_c471_6e5e_4fb4_ab31;
        state = 128'h0d0a_65a5_f312_ecc8_c757_79b5_c51d_cb0c;

        #200;
        key = 128'h59ae_7cdb_af67_b597_0a02_f780_fd55_4226;
        state = 128'h6595_e09d_720a_8354_5939_88f9_e360_292e;

        #200;
        key = 128'h9f47_95cc_b92c_3774_4edb_a09d_9a66_9f7e;
        state = 128'h5ba4_8ab7_915e_8de4_4d97_3e0d_b355_8d49;

        #200;
        key = 128'h44b3_68c0_8512_fcf7_8701_2a5d_a8bd_5e60;
        state = 128'hfbaa_c244_e7a7_2d59_9eba_4022_6436_e4ae;

        #200;
        key = 128'hefef_fa36_ccf4_9f8b_6d4a_c533_7761_c353;
        state = 128'hfe20_224c_aa3c_0859_b052_7dc8_dfb1_05e9;

        #200;
        key = 128'hcfd8_79dc_8242_116f_ea06_be9a_955e_96b6;
        state = 128'h5b0c_9e36_106e_252c_dcfa_cf2c_b05b_ca72;

        #200;
        key = 128'h3778_0410_105f_e9d8_3ed8_e321_42d6_1666;
        state = 128'h75e1_df99_7c02_156d_4e6b_a5e9_c742_3b54;

        #200;
        key = 128'h3df3_996b_1713_e4e2_a4d0_af40_e42f_567b;
        state = 128'hcbbd_158d_f636_f72f_839c_efc1_a029_00bf;

        #200;
        key = 128'h562c_b260_f055_f9d3_d0d1_69cc_d5c9_44a6;
        state = 128'h68fe_da91_8469_0a31_72b9_cabc_465d_969b;

        #200;
        key = 128'he856_48d7_ff1e_fc31_7587_4895_a4dd_8fe6;
        state = 128'hd4a8_e3c5_6636_8d1c_740b_47ae_000a_b712;

        #200;
        key = 128'he18d_6c43_c57d_4ab8_0829_b1c4_4cf2_32b7;
        state = 128'h33ad_3813_86e6_f033_3119_b2e0_00c5_1f45;

        #200;
        key = 128'h77ee_2893_60c4_653f_08b1_b05b_072a_de01;
        state = 128'h7b14_e746_c154_1753_8b4f_e508_449b_ce9e;

        #200;
        key = 128'h8181_2dee_6194_f223_8138_32b4_d14f_b0ca;
        state = 128'h86aa_2fd6_6eae_69f3_4be2_dc92_bcb3_cd74;

        #200;
        key = 128'h1790_a003_e333_d6de_996f_dcca_680d_b89c;
        state = 128'h3edb_951c_08a5_4ca7_39fc_3072_33e9_6b67;

        #200;
        key = 128'h98f4_d2ac_8bfd_1ef0_6656_bd5f_dfbf_9d3f;
        state = 128'hadce_3603_2928_e57c_23e8_7167_8a19_47ce;

        #200;
        key = 128'hb2b6_c9ad_b46b_17fc_574c_bebe_befb_1365;
        state = 128'h2d97_0fa8_acfc_bc2d_ef66_11ee_fda0_523e;

        #200;
        key = 128'he784_393d_ed6e_3e65_51ce_b712_cda3_c881;
        state = 128'hd3ac_d9eb_4c53_e16d_6b7a_18be_ca36_6fde;

        #200;
        key = 128'h0028_46e9_9959_27b3_d70a_ab34_9324_6888;
        state = 128'h3b6d_c503_00de_f773_316d_8347_c356_ca78;

        #200;
        key = 128'hc844_ba4c_327f_4c74_1214_a102_1a00_09d2;
        state = 128'h7be1_f475_f074_dc88_8a69_e49c_2ea0_7679;

        #200;
        key = 128'h1995_cf67_2dd7_99e4_e3dc_6f8f_fbc8_849e;
        state = 128'h4e15_7bfb_e09e_ee6e_4a74_bb37_f2c3_6387;

        #200;
        key = 128'ha8b0_b0a0_560c_4782_d010_5e72_816c_28e9;
        state = 128'hbd9e_17d0_e7bf_5b5a_efa6_1f83_ca68_de0c;

        #200;
        key = 128'h5e9b_e549_1f74_c3ef_e0ca_b9d3_4d57_2f47;
        state = 128'h2c9d_afea_b57e_13c3_f9a4_1fb4_1155_29a8;

        #200;
        key = 128'h6d83_37ec_2729_fa2f_a9e9_858a_ac85_c4ee;
        state = 128'ha2fa_ed88_7015_864d_957a_2714_9e9e_4b26;

        #200;
        key = 128'h3e82_8b63_73e0_4cd2_1907_6ea9_eac7_c72a;
        state = 128'h6211_e4e6_125a_8d92_6dd7_71b3_cde4_1635;

        #200;
        key = 128'hbb6e_60ae_f830_7c9d_233f_793b_6cad_1f3e;
        state = 128'hf422_fcd8_c876_ee83_9f35_9e07_d13a_0b6b;

        #200;
        key = 128'h9719_7b12_0bb0_6c89_cb67_8d4b_1b48_cb46;
        state = 128'h32ea_57e4_2f2c_83fd_d341_c137_e683_4240;

        #200;
        key = 128'h11b2_9d46_fdab_9c99_528d_2067_f923_7663;
        state = 128'hf6b9_72be_8c8d_f3cf_e576_2c3d_7eab_1c9b;

        #200;
        key = 128'h048f_f696_9961_b553_1e25_c615_0c5f_55ef;
        state = 128'h11c7_0830_1eb5_eb28_2f95_a86a_e76b_8dfa;

        #200;
        key = 128'h0e3a_28d4_c037_fb59_9bbd_9ae3_ef4c_5571;
        state = 128'h6e80_de73_3b65_e23b_1dca_a6fa_daf3_cc54;

        #200;
        key = 128'h49ff_9cdf_4182_f189_dcb7_918c_083a_b654;
        state = 128'h268a_e754_9490_739a_d582_7e88_9480_c904;

        #200;
        key = 128'hc255_ec34_a06b_8eee_f88a_e3aa_f8b5_85fe;
        state = 128'hc880_48ab_deac_f112_895e_b6d7_c540_5201;

        #200;
        key = 128'h21c5_4c1d_cba2_db67_a99c_7bd9_eec8_7c69;
        state = 128'ha1bd_f992_595e_2f50_a6e6_bef4_a8dd_b450;

        #200;
        key = 128'h28f8_c930_2763_35f8_8ec3_98a8_d398_563e;
        state = 128'hd7d0_968d_0386_d766_236d_0a62_4152_44e7;

        #200;
        key = 128'h22f6_ab61_b440_948f_13c3_e5c6_15c7_47a8;
        state = 128'hd651_edaa_ce13_7ed5_d6fa_9dd6_aae8_099c;

        #200;
        key = 128'h53f9_86de_2113_28ca_2832_2c29_0642_1360;
        state = 128'h694f_98ba_271a_3a8a_d610_bcf4_c478_3d9a;

        #200;
        key = 128'h3b0c_90f9_f86d_d8ce_1c6f_b835_496d_1eaf;
        state = 128'h03a9_6667_2fee_2280_f6d6_1305_7ae0_d1a0;

        #200;
        key = 128'hd4c0_f61a_b4de_9adf_9247_88fe_2630_d8ce;
        state = 128'h3841_25c5_ab34_52b4_82f2_918d_0898_5106;

        #200;
        key = 128'h4caa_3994_805d_3a88_7de0_b28e_d3a8_ac31;
        state = 128'h2805_0d0d_736d_f607_7753_84f1_f111_0522;

        #200;
        key = 128'h731b_4485_84e1_09ea_2d1d_460b_d095_7f61;
        state = 128'h048e_2a27_2300_111b_57fe_8bc7_56d4_b869;

        #200;
        key = 128'h6fb4_eb90_135f_5886_df57_b4cd_a61e_29ba;
        state = 128'hfb1d_2db9_372d_04e6_b5d0_7049_da7f_6bb0;

        #200;
        key = 128'hfc1e_dcff_10c5_4628_d306_419f_561a_f025;
        state = 128'he977_d1bd_fdb1_0512_3584_5885_0899_437e;

        #200;
        key = 128'h6efa_b416_7ea8_00c0_c36b_7e2f_046f_0f93;
        state = 128'he62e_9cc0_c4b9_ca99_273b_e8e7_0d59_b678;

        #200;
        key = 128'hd171_1234_66d6_e759_f9ac_53dc_2d93_f221;
        state = 128'hbdca_8a30_36cb_7cbb_e5bb_6fad_54ae_fe84;

        #200;
        key = 128'h5970_2a7b_6766_043f_65cb_3f75_4a14_05c8;
        state = 128'hfe5f_cada_a2c2_ba50_5628_1af3_d9ed_0d46;

        #200;
        key = 128'h7a72_5990_f861_01ef_f94d_0c24_cbcf_f69f;
        state = 128'hcb3b_3731_a2a2_12a3_ead6_5d9c_29bc_15c6;

        #200;
        key = 128'h17b5_3242_5ac9_c09c_2b72_b670_41e1_bb74;
        state = 128'h57c7_ba69_ae38_099b_5e34_9115_58b3_30d9;

        #200;
        key = 128'h3f26_ae40_e1b4_d75c_97e9_b601_e543_0690;
        state = 128'h1ed2_d469_bbcf_9e06_604d_f962_deca_f9a3;

        #200;
        key = 128'h1186_797a_2635_c2ec_21a9_b669_05b8_439c;
        state = 128'h14a2_5c24_9343_d7f1_ea6d_9533_ec49_bfe8;

        #200;
        key = 128'h1b18_7f0a_feed_e4e4_1db8_b74e_b952_2e5a;
        state = 128'h610a_0355_5fc5_8228_f36f_6778_ad5b_a0ea;

        #200;
        key = 128'hc9f6_c14a_0ff3_7f51_9666_5340_954d_dbcd;
        state = 128'h9a8c_7313_7e4c_c958_a901_d5e4_ab74_e2dd;

        #200;
        key = 128'h20f1_ade4_58f4_e623_7997_6fb9_a135_35c0;
        state = 128'h5cf1_34c8_d5d3_a880_7a71_04e5_6d4b_59f5;

        #200;
        key = 128'hf3f2_779e_fb0d_1e5c_9f7a_07d4_fbb4_fe5a;
        state = 128'hb912_c0c5_5277_4ad9_a39d_8d4f_2961_12b5;

        #200;
        key = 128'hc602_ccce_eefa_a7b2_c64b_ebf0_566a_6745;
        state = 128'he81d_1efb_9eb4_9916_4757_ce98_436e_c2a7;

        #200;
        key = 128'had8f_c1ed_2af5_6470_9956_9521_5ed7_914c;
        state = 128'hceeb_ecf6_a2fe_fb8a_c571_7be0_7545_f4c0;

        #200;
        key = 128'h4e60_e925_d06e_704d_e99b_3a17_ecd0_98c5;
        state = 128'h13dd_ebe0_af32_2aa6_1ec6_7c09_fc09_4a52;

        #200;
        key = 128'hf302_9e70_ab2e_049a_c203_17e6_6cf5_3791;
        state = 128'hea91_3542_e8a5_a8ea_1050_255e_870e_0684;

        #200;
        key = 128'ha5e9_77c5_de58_b74a_3dcf_ff3e_fa63_ef33;
        state = 128'hdeb6_e976_282f_9e2c_8f03_8c1c_8919_2fd3;

        #200;
        key = 128'h7163_9dcc_3544_29b9_b76c_e7e7_26c4_dd8b;
        state = 128'hfbf4_3445_0b4f_f385_1519_f211_b2f2_156f;

        #200;
        key = 128'h7e9b_7355_dd8e_3e4e_15bd_0456_bf1d_8ce1;
        state = 128'h820a_c3e9_cf5a_e315_213d_3ffb_9aec_d66c;

        #200;
        key = 128'hffcb_b70d_a509_691d_e494_0bca_8cab_2ec6;
        state = 128'h0099_d47e_0002_b9c4_c7c1_4582_a4bd_21e9;

        #200;
        key = 128'ha912_5549_97f1_0ab8_e076_b8ca_a276_8c6f;
        state = 128'h1f71_fdbb_c894_fef9_1a0b_bf19_3615_16a8;

        #200;
        key = 128'h89e9_d956_9234_0fe3_8e70_5419_7882_4e61;
        state = 128'h474b_a792_90a4_53d5_36c9_b40b_bf26_cf5c;

        #200;
        key = 128'hc50c_19ee_8245_dea1_2b53_b226_53e5_ddc7;
        state = 128'h148f_cdd4_71e5_b2e0_fccd_540e_e941_0fa6;

        #200;
        key = 128'hf2c4_5861_6213_ec7b_d978_fa35_1eb5_7122;
        state = 128'h345d_3de0_2a94_ff16_9cfb_580e_5338_5fd4;

        #200;
        key = 128'h9055_784c_fa56_7f56_bf89_9140_67ee_884b;
        state = 128'h30d1_bb99_0b22_ac8d_bbc7_748b_c180_e23d;

        #200;
        key = 128'h056a_42cd_48b4_dc95_278f_5887_6595_880a;
        state = 128'hf6c4_aeaf_4cda_61f5_3a86_516f_1e09_75b2;

        #200;
        key = 128'hb4ec_90f0_e606_250f_2535_5ca0_4317_f4a8;
        state = 128'h673f_42aa_f77b_7be8_8789_4a8f_3520_dd1e;

        #200;
        key = 128'h9726_2dbf_ce78_30a7_b244_f664_b4ed_e891;
        state = 128'hfd7f_b95c_c9a2_2e7e_cff9_a1a4_b6f6_afc5;

        #200;
        key = 128'h1775_811b_d60b_a937_f978_b850_90d3_8f95;
        state = 128'h7442_f8a5_8da7_abb2_0606_e18c_7cc3_1259;

        #200;
        key = 128'ha4f3_45e6_8cf8_ce9c_1d9f_20dd_9c61_ec4f;
        state = 128'hcb6a_8a7d_e87c_e4f8_9245_51aa_284d_d72b;

        #200;
        key = 128'h11c7_21f8_26c3_3ce3_72c6_6057_0f02_0354;
        state = 128'h2024_66f6_0987_c5d6_1cf4_72f0_f1b2_42b7;

        #200;
        key = 128'h9130_7d31_f3ea_cbef_f890_422c_f8d9_2646;
        state = 128'hd7e8_374c_6ae3_6475_d457_805e_08c9_b33f;

        #200;
        key = 128'hb872_a5c7_77ea_251b_a995_7034_f9a6_c115;
        state = 128'h94c3_1537_3d3b_db8d_8e85_4d6f_97b3_1621;

        #200;
        key = 128'h48cf_3b0b_078a_679c_7b67_03ef_f79e_96aa;
        state = 128'hff22_0b1f_e890_74dd_0325_8629_dd43_e60c;

        #200;
        key = 128'h0783_ade6_3dfb_cb0f_c22c_b0d3_f7d4_ed5f;
        state = 128'h4e3d_b908_4a93_0f65_30a9_a4e1_d140_0745;

        #200;
        key = 128'h227d_8a6d_13ca_48ef_82ad_e64e_e4d3_a26f;
        state = 128'h0db7_f09e_769f_843c_d105_ad3a_8364_a668;

        #200;
        key = 128'h1ca5_692b_97a3_8545_02ea_9d60_b091_20d8;
        state = 128'hceab_4d4d_1ef6_ec9c_47ff_1a42_9278_6166;

        #200;
        key = 128'haa92_2ec1_4ea8_9e37_40dc_c2f8_df85_2e85;
        state = 128'h624f_16dd_cbaf_7ba7_2003_db30_d9b0_d78b;

        #200;
        key = 128'h9f42_6c39_8e9a_0f76_05e9_332c_73b4_9aab;
        state = 128'h0dcf_a51e_a25d_8fed_965f_7bbf_9e1e_46f5;

        #200;
        key = 128'h0bfd_7afc_e619_1973_e642_fc84_49d5_74c9;
        state = 128'h85f0_3a8e_19b0_6cc3_8b11_906c_4587_355d;

        #200;
        key = 128'h9a96_90e8_067b_ce0d_f0b7_cd03_755c_6fd1;
        state = 128'h0388_a7ed_2469_6eb4_4964_0a60_a6c4_100c;

        #200;
        key = 128'hfd30_e9d7_f98d_1d95_b359_bd22_a330_7b0b;
        state = 128'h24cc_33c9_3444_703d_cf7b_5895_b070_f659;

        #200;
        key = 128'h9b0f_9100_b049_f89a_f8ab_4a6a_1194_404f;
        state = 128'ha8af_7937_0956_ac8e_173b_5cdd_1672_371b;

        #200;
        key = 128'h204b_f13d_8ec4_2d23_5be1_d3cb_c71f_e8e2;
        state = 128'h7f94_20c5_8766_c3fc_3cb9_eb1f_6a11_1113;

        #200;
        key = 128'h75ca_4e27_fb7e_848b_3737_e6c5_90fb_aa5f;
        state = 128'h03f1_4fcf_8e5a_afb4_a8c7_ce72_4204_35a0;

        #200;
        key = 128'h3530_845b_fbc0_0e82_0ec9_2c21_6e98_7cea;
        state = 128'h461f_4cfa_bf09_25db_71a1_365f_cf87_9e71;

        #200;
        key = 128'h1563_f404_eea7_b982_3b33_3ff3_ab11_418a;
        state = 128'hf2e2_164f_917e_c611_feab_55e0_e396_d9ce;

        #200;
        key = 128'he10f_c2c4_68c7_11b5_ed68_da08_d684_9285;
        state = 128'h91f4_cb6d_1432_a14a_2de5_fbe5_88b5_8a75;

        #200;
        key = 128'hd0a4_b79e_d6f4_8c25_3dd5_f581_d96c_6d56;
        state = 128'h169a_3d80_cfd8_7df3_b663_20f2_2c94_29ad;

        #200;
        key = 128'h229c_011d_899c_ed43_088c_a1e9_6370_3bc4;
        state = 128'h3b58_7650_ad22_a962_4370_d5db_e761_791c;

        #200;
        key = 128'h4609_32cc_cf94_419f_f284_ab7e_3827_1d34;
        state = 128'had4d_d2b0_8068_83e5_b114_28b8_dbef_fa3e;

        #200;
        key = 128'hf286_98aa_f1ac_1172_8a5a_ae7d_d1a1_7fbe;
        state = 128'hfc46_d261_b2fd_15e1_8e30_6840_d61c_36da;

        #200;
        key = 128'h065f_d33e_8395_297a_3d7e_a67f_5a9e_71e1;
        state = 128'h6876_ac80_d3c8_c05a_ca16_fcd9_7d56_ab99;

        #200;
        key = 128'h0fe1_cbf9_30e5_93da_4d66_c193_3b63_dab7;
        state = 128'hd362_4576_68ef_ed93_4e99_1c3e_5c87_7978;

        #200;
        key = 128'h8fcf_cce6_2c73_8e36_0861_664e_e38e_f9ab;
        state = 128'hd4b4_73f2_6e42_d64d_684a_9a4c_d8e4_a7c1;

        #200;
        key = 128'h743a_7b26_c350_956d_7826_28a5_b2c7_63bc;
        state = 128'h6edd_cc95_4388_9283_5fb7_4b61_173d_1044;

        #200;
        key = 128'h2dee_8db3_e2aa_ed67_0ca5_49c7_2f0e_81e6;
        state = 128'hc567_c73b_e19e_3779_f98b_f9cf_1a84_51d3;

        #200;
        key = 128'h74b2_b130_fe24_dc40_8599_9a34_e9e7_e3c7;
        state = 128'h8562_4797_39f9_c1cc_177c_9213_1052_6db1;

        #200;
        key = 128'hff56_3352_b6af_9b21_0c8a_e4f0_fc51_da2b;
        state = 128'h9c24_2bcb_5ade_dce9_4cf7_c63e_7147_6d1e;

        #200;
        key = 128'h2e43_241f_de5b_49f8_f08c_e084_d3a2_84db;
        state = 128'h3b71_7ac5_ccd9_49d1_99fc_cd94_af16_8208;

        #200;
        key = 128'h26d3_df11_496a_659e_bdc0_98a1_8b4d_ea45;
        state = 128'hf2c7_5cf4_ec42_ee46_5642_e9b1_49f1_2fa9;

        #200;
        key = 128'h3741_1242_b400_8163_25a4_56ac_9eeb_eb70;
        state = 128'h8590_d687_427b_fdb3_4048_7998_2967_210a;

        #200;
        key = 128'hd563_e089_d303_88bd_10a6_e188_b356_4fac;
        state = 128'hda72_b683_17eb_9ef8_a3a3_e6fa_27a4_8d2d;

        #200;
        key = 128'h1789_ac0d_8342_bed8_8c05_d8a9_4f5d_3067;
        state = 128'h55d8_6d43_2715_0239_7ccc_65c9_8fbb_8cdf;

        #200;
        key = 128'h1033_a00f_3f5f_65b8_6f1e_b885_b3ba_385e;
        state = 128'ha97a_75e8_6e5e_a8da_a24d_8011_fc7f_7e81;

        #200;
        key = 128'h12d2_7683_1435_ae88_8b0e_6053_fea4_e25f;
        state = 128'hf14a_529e_36b1_fce3_64e9_0366_3b9c_8971;

        #200;
        key = 128'h005e_14c7_f857_6063_7aa9_120e_d366_5761;
        state = 128'h1744_d3a5_5263_90d4_d1cf_6f75_cc27_48da;

        #200;
        key = 128'h5559_e454_03cf_dcf4_435e_4272_59b5_24b8;
        state = 128'ha389_4460_bcd3_ebf0_c90f_d9a8_e9ea_a71b;

        #200;
        key = 128'h6d70_408f_4605_c9df_b048_c8b3_4b78_0e1b;
        state = 128'hefeb_d721_da88_9f5f_beef_a0ea_5110_d3f5;

        #200;
        key = 128'h158f_43e2_4175_1e96_890e_0358_3614_1ef9;
        state = 128'h68f2_cd67_ca34_ce5f_e019_62df_b930_00fa;

        #200;
        key = 128'h6e09_8ac6_637d_b4d5_2311_65da_7fe3_55eb;
        state = 128'h74a8_a7f6_4c48_4698_cadb_7fe0_0b7d_2a3a;

        #200;
        key = 128'hcb43_38c1_0ef2_dd32_c2c0_6008_196d_7c57;
        state = 128'hbdb2_e97b_725f_88ce_e5ca_0a37_ad9d_d36b;

        #200;
        key = 128'h72f1_d6ec_f259_ad9d_6dc1_db10_625d_01f5;
        state = 128'h6487_530c_e265_5935_a98e_f236_3a53_87ab;

        #200;
        key = 128'h9efa_c6e6_c932_38a4_f14b_d282_ecd4_1f04;
        state = 128'h9af5_bb4e_8653_55f1_e727_dc0c_c086_e92b;

        #200;
        key = 128'h5574_dbf4_c004_41bf_2072_045c_b177_d74f;
        state = 128'hf332_2081_a968_86c1_8a77_eac9_55c7_e5f2;

        #200;
        key = 128'hdcf6_edfe_8b21_145e_eca9_00a9_26d5_6cc1;
        state = 128'h65bb_be98_b0f0_dd64_08d6_4c77_4cd6_141f;

        #200;
        key = 128'h9caf_d2d6_f601_0787_74a0_67c5_6123_4ae4;
        state = 128'h4b17_ffe3_baad_e916_aa26_0de0_a1b7_f50f;

        #200;
        key = 128'h6c7a_1709_07e5_e325_cbf3_3549_951e_a5ac;
        state = 128'hd273_2ea0_241a_1249_e257_6874_ebd2_57c3;

        #200;
        key = 128'h1409_43a9_edf2_96f3_66fd_c436_36d2_0d2e;
        state = 128'hc1ed_f8b0_555b_6e4e_8899_096a_b568_4624;

        #200;
        key = 128'h69bf_b463_4fc7_d98b_d6b6_e5c3_8d05_f200;
        state = 128'hc94b_2745_9b35_b831_0eec_9117_c88b_781c;

        #200;
        key = 128'h6c17_b0a9_765b_b523_4bc9_c0c3_5b81_1c6a;
        state = 128'h458b_878c_0b32_6422_bf91_5714_777c_d045;

        #200;
        key = 128'h2517_4126_e33d_03c9_4cf4_1c82_03b3_f03f;
        state = 128'h846a_36b0_4ccf_38d0_9138_537f_14a7_f22b;

        #200;
        key = 128'h41a9_5f87_bbec_9241_ec2a_7738_924b_8c33;
        state = 128'h81d9_1f23_42fc_527e_4d5a_14dc_4294_4735;

        #200;
        key = 128'hb223_a473_2842_7798_8283_e85f_3968_0ca2;
        state = 128'h2e18_9f2a_61b1_be07_6566_fadd_ea62_85a2;

        #200;
        key = 128'h0481_3181_31f4_f558_76cc_b085_0ad0_5833;
        state = 128'haac1_aad7_3cda_bf81_6f86_7ffa_1e51_8197;

        #200;
        key = 128'h2f54_305e_b6f1_02ee_c08d_6b55_5c5e_1e7d;
        state = 128'hb981_b7b9_5257_3f6e_5c11_138e_da43_9b21;

        #200;
        key = 128'h9e5a_0a57_c675_f0d5_4d01_5c75_dbe2_5e8f;
        state = 128'hb81d_8277_8abf_4c66_b2dc_fe67_8d82_be09;

        #200;
        key = 128'h2ac4_e715_96a0_1ed8_3a12_4d3c_a8fc_00aa;
        state = 128'h240b_f4f4_355b_f670_47bc_6c63_37b7_dc06;

        #200;
        key = 128'h92cd_2069_d68d_9efb_c972_2201_a791_f9fa;
        state = 128'hc9d4_9b07_2b9f_c972_cb54_120d_839b_6561;

        #200;
        key = 128'h0438_cec5_7c6b_8d23_6508_9d9f_7c34_555d;
        state = 128'h404b_e47e_d8c3_85fc_d2fe_038c_ccac_2cb1;

        #200;
        key = 128'h7989_1462_eddd_d34d_4cf1_eef6_c1ae_380f;
        state = 128'hd114_b908_b58a_390a_763b_582c_399d_996f;

        #200;
        key = 128'h34cc_3f75_3516_3f6e_8eae_3124_f9be_3fa4;
        state = 128'hac51_c6c1_653b_4fe5_a212_8743_5ab3_cf4b;

        #200;
        key = 128'h10a0_bfd3_532e_bdfe_53ee_21d2_ccb0_e3f2;
        state = 128'h8374_a4ae_2865_cfb5_4b1e_ac13_7102_afff;

        #200;
        key = 128'h29e7_7101_2b7f_3f4f_8acd_28c6_08dc_e1dd;
        state = 128'haa95_c5c0_e4b1_3ab3_06db_7149_78f6_ad68;

        #200;
        key = 128'hdcc6_1bdb_a3c9_1400_e227_6aea_f5cc_b84f;
        state = 128'h7989_48a7_7e2a_c5b5_1cc9_9247_c061_038a;

        #200;
        key = 128'h26a9_e363_be16_0bf0_3047_f439_8f97_75cf;
        state = 128'h8c57_0438_ac88_12ae_5249_f163_d3dc_1e6a;

        #200;
        key = 128'hf7cc_f57e_4a1a_56b0_ea94_6625_26d9_efc7;
        state = 128'h88d5_80e8_725e_63cf_ba6e_1391_863e_88fd;

        #200;
        key = 128'hbea0_b571_8630_b440_5c27_d2b5_c0d8_8834;
        state = 128'hfb73_8e39_dd06_134b_46e5_0837_cdfb_1c3c;

        #200;
        key = 128'h2a54_0426_4c5d_c2ef_80c9_ed57_208c_1f46;
        state = 128'h6ad5_ed0f_5c56_97f5_8192_5fe6_5993_db61;

        #200;
        key = 128'h2c94_9d0e_4d23_aa8b_828a_647c_8446_3fee;
        state = 128'h9c7b_2d09_4c7d_ebc7_0bfb_1e56_19e8_9033;

        #200;
        key = 128'hd47d_a3de_9e86_19cb_7dc4_4413_34cb_88c1;
        state = 128'h4a58_5af8_6cbc_add0_9c2c_bcd4_e92b_0880;

        #200;
        key = 128'h9380_e103_f378_7243_62a2_14cd_18fb_bdba;
        state = 128'h97e0_48d8_35c6_2dfd_f019_aa13_514c_ea81;

        #200;
        key = 128'h17fe_72e2_74a1_4e75_e515_2e85_1bfb_e210;
        state = 128'h41b4_2208_6db3_4c1a_60b8_f0b8_9cc1_e9af;

        #200;
        key = 128'h2934_0ef9_e96b_e178_91b2_d783_862a_a444;
        state = 128'h8229_bfa2_9115_c7ad_4bcc_8e07_8ab0_d944;

        #200;
        key = 128'h3dac_2eaa_f6fb_d1d4_8f87_1420_6341_53b6;
        state = 128'hb411_2b96_5ca1_b4f0_1344_514f_c63d_2e05;

        #200;
        key = 128'h52ef_5ff6_67fd_e5ae_d83d_2968_1b09_f972;
        state = 128'h8441_73f6_9a56_82ba_1eea_bbbb_7375_552f;

        #200;
        key = 128'hb939_1912_275f_834b_4449_13b0_f0e0_091d;
        state = 128'h6121_0089_5441_8cf9_f46a_6731_85f1_889a;

        #200;
        key = 128'h77bb_edda_b826_e918_98a6_69c8_295d_8d73;
        state = 128'hdd21_3a99_6855_ff4d_4877_4bd2_3e53_d028;

        #200;
        key = 128'h0e36_ba20_e8a2_0f37_54a4_6519_4554_be2d;
        state = 128'h3015_ea38_6e9a_80e6_7e0f_83a7_c401_738f;

        #200;
        key = 128'h03dd_d5fe_d2b1_ccb9_a2fc_2af2_2c4c_10a5;
        state = 128'h4ef8_7282_1307_3c96_20ff_2e15_075b_2b48;

        #200;
        key = 128'h233e_b33f_9d09_a217_5364_36e4_4689_8fb0;
        state = 128'h9f5d_e1b5_b8e4_d705_1ad2_f6de_e50a_694c;

        #200;
        key = 128'hd54b_8db4_fb32_d235_06cc_277d_1401_c8a1;
        state = 128'h8517_350a_4f7d_43ef_2702_76da_00b9_4e17;

        #200;
        key = 128'h858a_f185_defb_a9cc_2869_9483_4273_d073;
        state = 128'h6e84_2185_8d63_ddeb_6b3d_9d98_92be_04f2;

        #200;
        key = 128'h8c36_3fff_e790_407f_d3cb_f1ad_066f_d060;
        state = 128'h2d89_0f6a_d7ca_f168_2857_b97b_4e7e_907b;

        #200;
        key = 128'h31b6_e23b_8020_1654_7e77_a096_aee6_6bb0;
        state = 128'h6528_dd05_5c0f_6158_1f4b_4167_e5e7_d676;

        #200;
        key = 128'h3c4a_b346_5e0b_3706_4aa5_4b83_cd4a_7bdc;
        state = 128'h3131_8bf7_6f6a_f074_fef8_f600_8a96_3791;

        #200;
        key = 128'h51ff_a02d_ae4e_5522_a807_b4af_c4f7_95c2;
        state = 128'h9c79_a9e3_4aab_ffcf_50df_8f8f_81a1_5921;

        #200;
        key = 128'h0841_4572_33c2_f75e_63d6_dd19_ee23_09cb;
        state = 128'h5a4d_b2dc_2e15_32a7_9bee_f272_03c3_b5a4;

        #200;
        key = 128'h9256_c728_c7bf_818c_5851_d9d0_a2fc_603d;
        state = 128'h68aa_1f2a_f8b5_2437_ba63_fffd_0389_8951;

        #200;
        key = 128'hffdc_5053_c465_cc98_e691_b113_2084_7468;
        state = 128'hf467_5d6e_c894_fdff_cc16_862f_0c62_c43c;

        #200;
        key = 128'h3ba8_3697_8749_569b_55d7_8e6f_3548_f29d;
        state = 128'h597b_fb85_87d3_530b_b929_fa6d_d471_e66a;

        #200;
        key = 128'h02ea_fb55_61ff_33f3_cd95_2070_42d8_b216;
        state = 128'he3a9_9a9a_bd40_5683_5c6c_06c0_6b67_d247;

        #200;
        key = 128'h8df4_0e9e_29a0_1268_6d48_7716_b660_039d;
        state = 128'h0836_b16d_0466_3cb9_c88b_08af_5cbf_5ae2;

        #200;
        key = 128'he73a_0497_5806_395e_fcfc_7249_2495_22b2;
        state = 128'hf606_05bf_935c_f32f_864b_84e6_0a67_bd5a;

        #200;
        key = 128'h5758_6cb4_15aa_782e_c8b6_b31e_08c5_5494;
        state = 128'h8e2a_2116_a886_9041_c641_7d1c_a248_4baf;

        #200;
        key = 128'h82ce_c51b_b338_29d0_8cba_acd7_a24d_c6f1;
        state = 128'h30ef_0ebb_52fc_49f2_30eb_bd8f_af71_c185;

        #200;
        key = 128'he712_f337_a6dd_3cd9_933a_c6ef_0e0f_6469;
        state = 128'hc763_b7dc_6570_dd93_5c88_248f_6c60_c2c9;

        #200;
        key = 128'hbf7f_f1a6_fdd2_d356_1ad9_a7d8_8105_9307;
        state = 128'h8ed8_02d1_839d_a36d_ff63_6fa3_8e8d_2548;

        #200;
        key = 128'h2047_f684_e527_752a_c2dd_84a3_10af_0196;
        state = 128'h8b4c_3cd0_6f03_8660_3860_f853_f337_d882;

        #200;
        key = 128'h9618_0e91_7175_85e9_9af2_6d03_77a2_66db;
        state = 128'hef41_9f30_bfc7_ec2f_fd9a_cb46_f0d7_9cf4;

        #200;
        key = 128'h05fd_dcaf_6447_36db_c24f_6d98_2278_e45b;
        state = 128'h9841_da10_cf59_3934_8644_6f57_63d9_3f8e;

        #200;
        key = 128'h3354_a1ea_12cf_799c_41af_6259_c39d_c0bf;
        state = 128'h3961_5cb3_f80d_ddaf_d3a4_8808_ea61_c11a;

        #200;
        key = 128'hd3dd_689a_ca71_7a2f_0cdb_014e_2161_9942;
        state = 128'h5155_4028_0a7d_8a3b_7058_04e9_9346_52a0;

        #200;
        key = 128'h42cf_5e14_259f_cc9d_3176_2130_5896_b4aa;
        state = 128'ha57c_0f8e_827f_60b0_d3be_eb8a_c765_d940;

        #200;
        key = 128'h57ad_6f2a_c4e5_e3aa_21a4_6fee_f7c9_1ec3;
        state = 128'h3281_8929_a722_8525_35af_2e4e_30c4_b16f;

        #200;
        key = 128'h109d_edda_314a_5f09_dc1b_77f5_ae57_4de3;
        state = 128'hb735_bcdb_17cf_4495_4b71_ee05_a7e0_eb74;

        #200;
        key = 128'h16e9_71e3_913e_1eb9_5c86_809f_4a6d_ba87;
        state = 128'hd400_b2b5_06dc_1086_54f1_2d9f_2ed7_e7bd;

        #200;
        key = 128'h3f45_389d_1882_f46c_1685_7664_fae3_9177;
        state = 128'hf599_a040_213b_f061_b798_98cf_5297_5303;

        #200;
        key = 128'he531_06ac_8e35_02e7_4701_cd58_9c0e_6d5a;
        state = 128'h9722_ebbd_91c5_65a8_9e95_5c86_e4ab_f1b3;

        #200;
        key = 128'hdea0_c4a4_6759_3aab_0256_6328_f1ed_a913;
        state = 128'hd49d_3b3c_3927_3cf4_d760_176f_062e_0e5c;

        #200;
        key = 128'h6455_7305_3e4e_1a25_3ff9_819b_e7c6_b802;
        state = 128'h1d57_9a4c_4ea9_94c9_2f32_909b_104a_2ba4;

        #200;
        key = 128'h98b9_9565_aec7_3f1f_631b_266a_8ad7_3cc4;
        state = 128'ha97d_0295_bde9_e401_6d6b_9a70_d69b_0603;

        #200;
        key = 128'hf22e_c712_5b66_b3b8_c243_91b4_fe79_d99a;
        state = 128'h926e_805c_3028_e946_c7d8_6436_a0de_3721;

        #200;
        key = 128'h045c_563b_a05e_5145_dfe2_e0ff_5964_8d70;
        state = 128'hcf0a_bc3f_ba58_f9da_c916_986c_0087_453a;

        #200;
        key = 128'hee28_ddc7_8e50_53b4_9861_28c4_4028_9fd1;
        state = 128'h438b_5be1_9971_b36b_6543_74a6_e36f_fcce;

        #200;
        key = 128'h13ab_2ff3_6fc6_7b8e_ab0d_a3e7_f601_4838;
        state = 128'hd538_52ca_ca47_0740_160a_e192_bfe5_7b32;

        #200;
        key = 128'h43ee_adcb_9c12_22d0_d6cb_acd3_b15d_a334;
        state = 128'h0d34_578b_9c53_d7e5_a83c_d318_b2a2_dad3;

        #200;
        key = 128'hab33_2b55_1224_2ad8_69fb_58bc_1a19_d056;
        state = 128'h1527_96f5_5da3_0766_2f51_4d30_9a77_b291;

        #200;
        key = 128'h224b_c967_8cc5_e763_19f9_795f_1da6_96d6;
        state = 128'he971_4971_fd07_7bcb_01c2_aac2_5b7c_155f;

        #200;
        key = 128'h241a_594b_09a0_4e02_344f_7b62_dc64_2903;
        state = 128'hf913_82d2_d0a5_4235_fe6d_7be5_87e6_7a95;

        #200;
        key = 128'h818e_7416_9d9d_6f9f_42db_2f29_d8d6_2e6f;
        state = 128'h3e2c_8cb6_819b_2847_0b07_0d44_879a_4f22;

        #200;
        key = 128'h0779_c4d0_4a96_f7f2_5cc1_fd96_3682_00e8;
        state = 128'hf191_d2d8_913f_441b_4c52_1362_6719_3e79;

        #200;
        key = 128'h00e6_e6e6_cf6d_a21b_40be_898d_8927_fe5e;
        state = 128'hc580_a872_684e_e3ed_ec7d_9bc2_3931_51b1;

        #200;
        key = 128'hc761_b74d_42da_18c8_c1d1_def2_92e1_3244;
        state = 128'hda0f_2fbf_2e5d_a603_8b50_c691_ba2e_8707;

        #200;
        key = 128'hbc76_be11_7367_0df6_6f52_3d0f_80a1_339b;
        state = 128'hd696_ddc5_1442_f211_06d3_0a03_c863_3b9b;

        #200;
        key = 128'h652d_1427_6d11_a600_6161_b840_658d_9398;
        state = 128'ha600_6c78_bc58_b95a_5ce6_5c46_a788_bed8;

        #200;
        key = 128'hd908_2b50_4e10_d942_26b9_f2d3_81ce_7ad4;
        state = 128'h1ed7_42f4_c90c_e5c2_9517_62f1_856b_20ea;

        #200;
        key = 128'hfa1b_40c1_05da_3866_a828_ebb8_b146_f67e;
        state = 128'h48f6_9437_f0f1_2927_dc5f_c388_f851_34e5;

        #200;
        key = 128'h247a_37ee_597a_e2a5_0ce8_6c61_0151_77fa;
        state = 128'h09cc_2195_c731_afb7_29e0_23c7_5fe7_3ef9;

        #200;
        key = 128'he6df_b753_d264_def4_eb70_c47c_0c90_ae41;
        state = 128'h45bc_0f2d_15b8_2aa8_c6f2_cc6e_31ee_ea7d;

        #200;
        key = 128'hba68_8270_cc98_67d1_f2f7_799e_6c24_ac87;
        state = 128'h98db_efc6_30e5_cab7_caa0_b126_8ae1_19ef;

        #200;
        key = 128'h6701_2c99_9f8b_cdf1_7dcd_7c62_fa5a_fd8a;
        state = 128'h580b_d2b6_c1f4_b24f_3a24_e3a2_d941_8db7;

        #200;
        key = 128'hde01_8dca_04ed_79b9_8751_343f_db94_5c8f;
        state = 128'ha3af_fa1e_831f_0725_b583_8ed0_e4e0_fbf4;

        #200;
        key = 128'ha6a6_7b34_92da_dac0_2f8d_c8d9_37cc_0898;
        state = 128'h1c99_1737_76d9_ee25_bb2d_836b_0caf_cae5;

        #200;
        key = 128'h30bb_dfeb_095d_8990_5594_9076_6148_c3b2;
        state = 128'h0bce_39b8_0e5d_7fb4_e997_04ed_4c08_73bb;

        #200;
        key = 128'hd386_5208_1bd1_0afb_0693_7221_4e53_2b7f;
        state = 128'h7886_9b46_7887_87b7_b77e_9c40_02a3_4e7b;

        #200;
        key = 128'h2e55_68cc_6345_ddd8_f176_0620_1c15_0cdc;
        state = 128'h10d9_c572_61b0_3c91_80c7_9613_999a_6d39;

        #200;
        key = 128'hdf7c_0203_ced4_513f_65a1_0344_2f61_bad6;
        state = 128'he540_cd35_5af3_6783_f344_1709_4c72_3b43;

        #200;
        key = 128'h5965_7e2f_6039_6fed_fb9a_f19c_36ae_1a23;
        state = 128'ha8f5_3a00_1f08_2613_51e7_8bf6_0665_b4e2;

        #200;
        key = 128'h51d0_4d73_84fc_7c02_9e9e_d045_595e_0382;
        state = 128'hf03b_2640_c3a2_811d_5f82_015e_f995_f9a8;

        #200;
        key = 128'hfb48_f5eb_1b71_d04e_67b2_696e_b40d_107a;
        state = 128'h356d_2397_ef13_26d6_23c0_bd5d_441b_bdf1;

        #200;
        key = 128'hb11e_fa50_a895_84bf_9583_276f_6b6e_3afc;
        state = 128'hd458_2563_d399_1903_4270_0cbc_0b11_782a;

        #200;
        key = 128'h3115_191d_b365_06c8_c1c3_2dab_ba9b_350e;
        state = 128'h1b33_1b95_20fb_db1a_7e99_18fb_db1d_216b;

        #200;
        key = 128'h9978_1a7d_8fab_9be4_bf92_cd8e_33fe_98be;
        state = 128'h52f5_d880_d8d1_440f_76e3_456c_bc4a_861f;

        #200;
        key = 128'h8a1f_1243_ebad_6ee4_733b_7765_dd64_988d;
        state = 128'h5531_3366_9dc8_2a76_87a2_ebbd_bd07_29fa;

        #200;
        key = 128'h608a_6970_a9c0_067b_d7f9_ea3b_d083_3f99;
        state = 128'h1512_b043_96aa_ff44_296a_e250_5220_525b;

        #200;
        key = 128'h9b6f_b281_d8dc_030f_f8a3_af54_f040_3ef1;
        state = 128'hd06a_78b7_f233_70ad_3e01_1637_92a5_73a5;

        #200;
        key = 128'h28d7_d6a7_7fdc_dea0_cc76_4515_44b9_221f;
        state = 128'h275b_372c_d2cf_349c_c2b9_1751_7f30_e602;

        #200;
        key = 128'h7edd_a4a2_e9e1_19b3_0e90_239c_e2ab_bd2f;
        state = 128'h47fd_a699_cd97_16c7_485d_507e_9c23_a5f0;

        #200;
        key = 128'h04f4_fbd6_7baa_3fa5_3877_eeba_67ba_6372;
        state = 128'hcf22_a269_3344_0ba3_2c47_8112_4df2_153c;

        #200;
        key = 128'h856b_bb23_a67d_c67b_62f1_1572_4104_d00e;
        state = 128'h332d_a94c_85ba_2a04_9692_5d38_37c4_bcca;

        #200;
        key = 128'h47f5_a465_5784_25b3_c4a1_06b6_9af4_e5dc;
        state = 128'hcedb_f59f_7466_fc40_2dfe_2862_692e_6b80;

        #200;
        key = 128'h4ea5_da5e_5eea_8eeb_c04c_7b79_1dae_0bc9;
        state = 128'hddb6_5958_24c3_7a81_cc69_81ce_d88d_2cfe;

        #200;
        key = 128'h5522_9281_c967_e119_b69e_37d9_3a5e_84b2;
        state = 128'h1d89_6a14_ba88_39c7_7d55_e614_4018_e489;

        #200;
        key = 128'h4a6b_7fe0_1b57_8f05_c3bc_c109_0b12_10c7;
        state = 128'h79f0_3ffe_7aba_cfd7_5c55_8c47_b1dd_ba5e;

        #200;
        key = 128'hf8e2_6628_67af_c1e2_ecff_0482_378e_cb9f;
        state = 128'h46aa_3643_78f1_22ce_5917_8898_346e_1d6b;

        #200;
        key = 128'hbb33_e01d_21f1_7cab_75dd_d53b_c4ee_9e2a;
        state = 128'hb67e_c1a8_e1b8_994d_63af_1649_0385_139a;

        #200;
        key = 128'hc54a_fb1c_09ec_896b_638c_a49e_649d_2e4c;
        state = 128'h7a8e_4426_1166_2dbe_2164_2d58_0c9f_aa82;

        #200;
        key = 128'hbd68_442e_43c3_185f_b608_b9c6_2148_2a0d;
        state = 128'ha497_b19f_ec80_57a4_6c91_2bb6_ca87_e9fd;

        #200;
        key = 128'h53ee_f00b_3597_422e_1fd8_98c9_4df2_eb3a;
        state = 128'hb09c_e8f8_828f_28c9_ffac_9585_ac62_4911;

        #200;
        key = 128'h74b0_fa92_1b57_6fe4_e3fe_c5da_96b9_4745;
        state = 128'hfb68_2f69_1706_81cb_b546_7381_2b2e_35c2;

        #200;
        key = 128'h1f71_a40f_ad3c_20b8_2017_112c_c868_8e1f;
        state = 128'h4087_2dd7_efcf_e49b_9b64_17c8_a955_392e;

        #200;
        key = 128'h6fda_c7d6_4392_14f9_21e6_5aec_4711_cb48;
        state = 128'h6be3_816c_ffa4_2d61_b0a6_4ab1_d243_0348;

        #200;
        key = 128'h8b92_b096_e7b0_4673_5dd3_64ed_9cb9_e60f;
        state = 128'hb1fd_b720_cfd4_aea1_0631_9d4b_8d48_6913;

        #200;
        key = 128'he2be_8f2e_c6cc_2d78_d751_22e5_672a_756a;
        state = 128'ha635_e21d_98f6_58f7_e4af_cddf_4c25_5948;

        #200;
        key = 128'hb36a_50e0_3f27_72a3_1cc6_25b3_22f9_542f;
        state = 128'h4f92_bc12_8f7b_9358_cdb2_8098_d6c0_0df3;

        #200;
        key = 128'h3906_6afb_20d7_06a7_3147_ee4c_057e_02fa;
        state = 128'h2cca_3fc4_2212_227b_0e6a_bd02_7cee_c0df;

        #200;
        key = 128'hd785_401d_dc1a_61d6_a855_ddf1_4822_cf74;
        state = 128'h7186_974e_473b_3f6b_202f_10bb_a53c_dc28;

        #200;
        key = 128'hcc0f_0faa_4eb7_941e_1134_c183_5176_4418;
        state = 128'h02ce_c532_704e_9c52_9e65_b782_b31d_fdfd;

        #200;
        key = 128'hc3ea_6e83_a33a_e2d0_2e87_cf0c_764d_5b10;
        state = 128'hf524_8894_5f59_e34e_7329_c876_00db_b1ce;

        #200;
        key = 128'hbf32_bb02_d833_cd2e_36c0_d660_f6a1_3209;
        state = 128'hb6b2_feaa_e88c_e9aa_9b02_c8e0_8071_39f5;

        #200;
        key = 128'h8675_1571_eaf8_d701_27e6_95ef_a9d8_de33;
        state = 128'h9da5_ce65_7305_2689_7be0_cd39_a1b3_28d6;

        #200;
        key = 128'h9845_f37f_8ede_0163_a501_bcdb_78ec_1a4d;
        state = 128'h62e2_b8e4_9d44_f0c1_2e48_bfb1_8cd1_4fe6;

        #200;
        key = 128'h9f71_badd_b8a4_8d96_2a06_7fde_748b_cda3;
        state = 128'h7d58_5f14_e403_0370_1e8c_6174_8068_6822;

        #200;
        key = 128'h10c5_9eea_6f87_3510_5cac_7c5e_fe0e_9007;
        state = 128'h96c8_7e45_921b_02d5_1149_e5fe_4db2_17dd;

        #200;
        key = 128'h5a7b_f658_04b4_95e7_c391_19c9_6082_d7bb;
        state = 128'hd6fe_4d13_3061_8c20_524f_2238_b2e8_c363;

        #200;
        key = 128'h36c3_7a7e_65b7_35f8_807c_711a_2ea8_5f83;
        state = 128'hc23e_ccba_c5f8_b5d6_9a4b_434a_99ca_ccaf;

        #200;
        key = 128'hc976_85c6_7a84_4bbf_0733_678f_f570_1d49;
        state = 128'h4b52_0db6_e0c2_4c3f_a1e3_144f_b465_e774;

        #200;
        key = 128'hc202_e604_6dba_f107_8783_69b7_410f_0b62;
        state = 128'h76fa_ad83_c581_857d_9d35_aa93_9ef4_5341;

        #200;
        key = 128'ha298_a393_5fcb_6860_e350_c3d7_0014_57ae;
        state = 128'hdfaf_e9d9_5f47_285e_2343_513b_7700_80bd;

        #200;
        key = 128'h30d0_13f8_efc1_3105_bca3_fb00_e115_500f;
        state = 128'h969d_401a_b975_6be1_810b_44de_01fa_dedf;

        #200;
        key = 128'h5d1a_ee54_284f_90ae_a695_3703_5f76_4296;
        state = 128'h751e_5b84_841c_6812_da01_aa1b_f9fe_2a5c;

        #200;
        key = 128'hbc54_0cc1_3af0_ef07_35ac_5b24_853e_0cfa;
        state = 128'haeb7_e6e0_ec0f_a7fd_0fad_3bdb_e309_dfa0;

        #200;
        key = 128'h7cc7_23fe_3d26_732d_8ac1_5ae7_1190_f542;
        state = 128'hc1b2_0ffc_90a6_937c_fe06_0d2e_5f20_064b;

        #200;
        key = 128'h38f4_f6b0_c014_0b67_6938_fe4b_3d91_e606;
        state = 128'hc421_2b6c_5d47_7033_a07a_09c7_64ce_6844;

        #200;
        key = 128'h7195_553f_a110_ddc9_1941_18b6_aee6_ea98;
        state = 128'h1834_abc0_7241_a19f_7ae8_0ede_77bf_6417;

        #200;
        key = 128'h1416_1074_1ab9_88a8_0f88_4aae_6f56_5e83;
        state = 128'h274d_85fa_82de_4a7f_a580_3f08_cddf_637b;

        #200;
        key = 128'h0154_912c_557c_9dac_23e6_5200_662a_803f;
        state = 128'h7268_5f65_8f5b_fff7_6066_e8c6_319e_51d5;

        #200;
        key = 128'h153e_512e_043f_3f5f_5528_c476_7cdb_8550;
        state = 128'hdf8f_5db9_b8c9_b224_8972_0a31_bdce_50a2;

        #200;
        key = 128'h7bbe_4e3f_2b79_822c_df76_2f8a_ee1d_0f27;
        state = 128'h56df_5ba2_16ff_c57d_8b5f_30df_c839_8b73;

        #200;
        key = 128'h4f73_fe27_c472_25ec_f2a9_f114_f6e5_ac72;
        state = 128'h1b5c_3fa5_53b4_a705_140b_f8d2_8e32_35e4;

        #200;
        key = 128'h85af_a0b1_16e2_af38_ab7d_86cf_d163_b274;
        state = 128'h8251_4101_aa98_991c_662e_41c9_f0d0_86ea;

        #200;
        key = 128'hd4b1_9993_4c6e_f947_11bb_37fa_c156_99b9;
        state = 128'h2b70_40ba_131a_6bd2_a31a_9a16_1703_7c6e;

        #200;
        key = 128'hc37d_bd3a_3f65_3e20_ff15_5034_7cf6_36f8;
        state = 128'h3585_51c9_afde_55d3_e57e_e570_da4d_c259;

        #200;
        key = 128'he4b8_497d_631c_3396_6c4b_7a44_e56e_d682;
        state = 128'h4b16_e64b_52f4_7010_03c2_d43e_c0ee_7db9;

        #200;
        key = 128'h24f8_abd5_4fc3_600e_7898_4080_4403_d6a9;
        state = 128'h6560_8bd0_deb9_5f5f_2ec8_ddfc_d54c_e997;

        #200;
        key = 128'h10ae_5cf7_b705_a267_c676_1321_aefa_9bdd;
        state = 128'h1578_34a5_8c1a_7731_4bc2_b2dc_f280_bd75;

        #200;
        key = 128'hedaf_928c_026c_760b_91c3_113e_83ed_f265;
        state = 128'h28b8_4224_de6c_72a8_229a_ed02_071b_4940;

        #200;
        key = 128'h96eb_9ab7_7bfe_d504_be56_dd9e_3381_12ca;
        state = 128'h77de_4d32_a168_01e4_d9cd_eae1_99e5_593f;

        #200;
        key = 128'h8c8b_ce1e_d027_ad31_6dbf_fcc5_eda5_d1b4;
        state = 128'h5fb3_ede0_c7f8_cdf5_8ccc_b7d3_8621_8a68;

        #200;
        key = 128'ha832_c5f9_b0e9_35b7_09af_6357_38b4_83fa;
        state = 128'h66b7_4282_48d5_88c2_ddee_cdb0_2881_c967;

        #200;
        key = 128'h5a2b_af99_868e_e588_c0ef_4097_1325_91ea;
        state = 128'habd1_38dc_5eec_7d9c_8c88_7a4d_ceb6_c95c;

        #200;
        key = 128'he2b6_f622_a3f5_487d_d707_1a56_872d_d639;
        state = 128'hdd88_774d_542d_2a1e_3621_6319_795b_0c15;

        #200;
        key = 128'h4f00_5f47_a8aa_f751_0386_aae2_3479_748f;
        state = 128'h74ac_5d3f_d7d7_1731_0212_d2cc_ed4b_5f15;

        #200;
        key = 128'hd1e7_52a6_db96_3db6_0a34_b716_6b94_e4cc;
        state = 128'hecc8_f4e5_2a12_8868_c38b_bd8d_8ee2_fb6b;

        #200;
        key = 128'h1d1e_e206_1f62_fd6f_1685_2ea8_094e_18ee;
        state = 128'h39e9_70fe_0e29_d355_dc39_b61a_fc04_445f;

        #200;
        key = 128'ha56e_8955_e19c_064c_60c0_9cb1_6e32_795d;
        state = 128'hdc82_936d_a1cc_5a93_e7d8_225a_213e_df12;

        #200;
        key = 128'h4e82_3adc_304c_91ae_2a18_0cf3_827b_0526;
        state = 128'h9d31_0e29_11f5_e429_a611_5103_0b94_8830;

        #200;
        key = 128'hb066_4ea4_aa15_3cc1_fdec_332f_be59_5998;
        state = 128'hc63a_6dad_2598_1e8f_3951_10ed_ed1c_ee6a;

        #200;
        key = 128'h94a0_cc03_c19d_63bc_8ca7_9183_b5fd_a072;
        state = 128'h0aa3_f824_c318_261b_b979_97f8_51c2_a2a0;

        #200;
        key = 128'h37fb_0003_6021_a263_eaa2_cc2e_0e72_16a4;
        state = 128'h248f_9a0b_17f7_c4dc_9a31_96c7_cf3e_8c7c;

        #200;
        key = 128'h6ab5_f090_e448_b09d_ff13_d840_9c66_f5ed;
        state = 128'h4905_625c_6661_d860_5a3e_3912_9b8a_db62;

        #200;
        key = 128'h3c68_b07f_3c93_5d6c_2cd5_7c71_79e5_b4ab;
        state = 128'hf569_4748_0af4_10ea_31ac_86d6_e7a2_c18a;

        #200;
        key = 128'hfa62_e057_8259_cab0_c2a2_f964_44cf_ca52;
        state = 128'h3b90_e1fe_1b69_8e8c_d9d7_242d_2a40_c789;

        #200;
        key = 128'hae7e_4759_5200_a157_b58f_218f_751a_022b;
        state = 128'h418c_0bf8_dd98_7966_2c4f_4822_3b0a_3066;

        #200;
        key = 128'hffc6_397e_9443_be47_e74b_4c60_ac3c_9ce9;
        state = 128'hd4f5_521f_1239_074d_cc4b_0563_8327_06a9;

        #200;
        key = 128'hedcd_d1f2_a8b8_0d97_1828_1acd_9428_0e2f;
        state = 128'h4a1f_68d2_e9cf_704f_d297_b93f_68de_914d;

        #200;
        key = 128'h0e1c_5b1e_6d77_98d2_fc5e_437f_44af_f853;
        state = 128'h8163_fbac_3ae7_86b0_6a65_2456_ea94_9431;

        #200;
        key = 128'hd2eb_bb3a_ec7c_89d6_6fe1_09ea_2de6_9b50;
        state = 128'hca69_6382_c574_2e99_dd18_1d54_8502_677d;

        #200;
        key = 128'h3f05_5dde_d273_f4ae_a04a_8cb0_3e65_83cf;
        state = 128'h9885_913e_c34c_8473_ea85_1111_4131_fee8;

        #200;
        key = 128'h4374_dedb_aa50_29ee_6fe0_5e30_1820_f425;
        state = 128'h5723_c33c_07ff_209f_c0b6_c216_363b_5b9c;

        #200;
        key = 128'he036_7bbc_53e8_9bbb_fbe0_48bf_2bb8_1938;
        state = 128'h54c3_5fe4_20f4_8115_963d_c299_db9d_7fbb;

        #200;
        key = 128'hf173_5d8a_850a_347e_2b83_a661_562a_603e;
        state = 128'h6333_6533_2f10_d4d9_6b79_66cb_248f_cc13;

        #200;
        key = 128'h8f52_0d14_9996_a46f_fe86_52f4_d411_340f;
        state = 128'h0943_6972_00b1_e91b_b14b_9df9_c569_5245;

        #200;
        key = 128'h0917_4826_c33d_0dd0_7cb7_3b4f_8dc3_f839;
        state = 128'h302b_a8c2_9303_9cf6_20f2_b31a_3f81_d779;

        #200;
        key = 128'h0534_cb08_3435_8b9b_b54c_7076_b87a_6932;
        state = 128'h9648_4e49_0427_dcd1_7750_2f3a_f7e7_6c57;

        #200;
        key = 128'h4906_3c65_bbf5_7096_ccda_594c_8f8f_3961;
        state = 128'h6735_b25e_6efa_58d3_9302_d26d_09a1_0db2;

        #200;
        key = 128'h8054_09f4_759a_0f69_cce4_0fb0_700e_ce11;
        state = 128'hd564_673e_bc71_c156_8fd5_66ed_b8a5_e146;

        #200;
        key = 128'h8366_77c9_9f3c_5799_66c1_3142_3b77_a8bb;
        state = 128'hda46_f1d2_2ea3_e825_c5f4_ce2c_110d_db75;

        #200;
        key = 128'h8407_55ae_fca7_b3b8_b085_74c6_c7f0_f4ef;
        state = 128'hd1bb_6f45_3ebc_113b_9527_4f36_b39e_38c5;

        #200;
        key = 128'h1479_bad5_72b6_6612_be8e_f0ce_caa3_06c8;
        state = 128'hdb85_a7f7_1c32_5724_1239_f8f5_2a5d_9113;

        #200;
        key = 128'h846a_e3b4_50f5_95e3_afac_bcb8_a757_c845;
        state = 128'h2f91_022b_8b71_3869_ea67_8f07_2c62_0c7a;

        #200;
        key = 128'h6846_9fa8_d31f_fa64_b7e4_1f7e_38e6_e9c8;
        state = 128'hc3d4_3371_344d_e68b_b83a_eaa9_6011_eb06;

        #200;
        key = 128'hbdac_6d45_31fa_d9ab_6a1a_fcbb_8113_9b4c;
        state = 128'h59bd_f899_72cf_6e88_61da_980e_bc04_1adb;

        #200;
        key = 128'ha5ff_c0b6_046b_7a6c_c261_d0a9_4fc4_d77f;
        state = 128'hc24c_8f9a_6841_4260_d553_1d84_1f04_4703;

        #200;
        key = 128'ha5ac_7843_acc9_1407_5ccc_f0f0_4942_da0a;
        state = 128'he234_a4aa_2741_7202_9495_a3d9_2bb1_f70c;

        #200;
        key = 128'h71cd_fb8a_2979_38e3_5e8e_9cc4_ad4e_a525;
        state = 128'h10e3_4267_b493_6e46_b3a7_9127_90a2_dba1;

        #200;
        key = 128'hc32d_4e9f_05ab_ee2f_7d25_8543_6466_21a1;
        state = 128'h45a7_4272_c7cd_0c2a_ff2f_3afa_0fe3_e403;

        #200;
        key = 128'h3262_0e59_2d7d_68b5_6988_a225_d615_ae99;
        state = 128'h0dea_29bd_2f6d_9d5f_6262_15e8_73d5_13d5;

        #200;
        key = 128'ha577_6878_849c_20ee_669b_39af_af59_2a9e;
        state = 128'ha266_95b6_ec4e_6360_c10d_aa5d_4d74_62aa;

        #200;
        key = 128'h2f37_1c43_517f_f42f_c68d_ab6d_2a8d_17b2;
        state = 128'h6799_c63f_2dd9_79dc_86e8_b04c_91ef_e68d;

        #200;
        key = 128'h95fc_3a55_1ffc_25f1_9607_47f2_7b31_35b1;
        state = 128'h2952_d203_ec16_6482_4217_9c49_6bd9_79c9;

        #200;
        key = 128'h3758_520b_2241_bc9c_b4c7_7140_7cd2_4291;
        state = 128'h73ce_6fcd_1c50_479c_b91e_da23_cddc_46c2;

        #200;
        key = 128'h86af_9579_15e9_a88d_b69c_46b2_42dc_4b1d;
        state = 128'h6b6a_b941_3cd6_d8dd_8f06_103f_c3b2_1297;

        #200;
        key = 128'h0b1d_454b_cdac_ca07_e57c_8db3_bf40_b989;
        state = 128'h1b57_c66a_e14f_1d66_d479_857e_e306_5703;

        #200;
        key = 128'hc015_fc14_1244_c9c7_7715_1b97_0ce7_b457;
        state = 128'hba26_2d77_ca27_58db_b77e_15b6_00bb_5960;

        #200;
        key = 128'h59b3_157c_6b89_21e3_ed70_cba3_47b0_2350;
        state = 128'ha686_7b32_e847_442e_d65c_bf47_e85e_8585;

        #200;
        key = 128'h8471_a7ac_1a1e_72d5_9f5b_2586_958b_b0ae;
        state = 128'hca5a_7edc_671e_b7d4_fe9c_73b6_82ed_81bf;

        #200;
        key = 128'he9bc_a56d_2115_66d1_5f54_bc0b_06f4_6ef4;
        state = 128'hd62b_de70_8fa5_02b4_1288_167a_7949_5c91;

        #200;
        key = 128'hf4da_9613_8651_c6b1_7807_c5e7_4abf_c5a3;
        state = 128'h1746_3491_c303_89a1_8a0b_f33d_aa7e_4a5e;

        #200;
        key = 128'hd33b_bd06_693b_48c9_447b_3d88_dec2_e52d;
        state = 128'h7c5a_ba42_5e7d_a9a0_85da_31e8_0268_a896;

        #200;
        key = 128'h9041_df23_b79d_67c8_6250_2aaf_2b18_eb8d;
        state = 128'h0daa_5029_df1e_a056_681f_dd5f_1529_e98c;

        #200;
        key = 128'he661_9ac2_154a_0e3d_271f_4910_2282_8d1b;
        state = 128'h7da8_7f2c_cd78_b50b_4346_f713_eb24_ce62;

        #200;
        key = 128'h661c_7340_cd40_5ff2_e54f_8051_d0e4_ab0f;
        state = 128'h688e_ba25_de81_c972_ac22_2657_3775_7d27;

        #200;
        key = 128'h1dbd_8003_db39_7b4a_5827_88aa_0f25_c85d;
        state = 128'h3f6b_49c2_ec86_9574_ce60_0114_46e1_2d22;

        #200;
        key = 128'hd5d0_6929_57a1_5782_6dd5_a590_e305_18bc;
        state = 128'h7ad1_1d47_1b56_8ace_2839_0b1d_3053_1eb0;

        #200;
        key = 128'h2dff_a18f_5208_ced4_0c21_2bc7_40e2_d417;
        state = 128'ha864_5fdb_91b6_e155_bb49_1fcb_2590_9b44;

        #200;
        key = 128'h0973_c92d_ac6b_4e67_d8b8_edea_e321_990b;
        state = 128'h8b76_9685_4f8d_54e7_038e_5c32_08de_e51b;

        #200;
        key = 128'h0ff7_3a10_217d_0430_7089_b854_7d24_6309;
        state = 128'h7e46_f6a9_af11_ccca_3f0f_afc3_b24f_3541;

        #200;
        key = 128'h4a3d_e031_a837_6686_8fae_684d_7bbb_1ff7;
        state = 128'h8678_26c2_e01b_5861_8a90_02f0_8cd4_c6ac;

        #200;
        key = 128'hb607_75bf_29cf_6724_aab4_3649_1a71_6039;
        state = 128'h57d6_23f8_8f8f_396f_1e43_aed1_e43a_78b2;

        #200;
        key = 128'hc2b6_ca56_31bb_5faf_3edf_375c_e6f7_e649;
        state = 128'hd162_cf91_aa37_6cc3_8cc1_e4ce_5eec_2b0d;

        #200;
        key = 128'h8ee8_77df_8e0e_80b5_ec9a_0ffb_7215_bc07;
        state = 128'hf699_ecff_4c0b_f9d6_5a21_4354_529a_6b14;

        #200;
        key = 128'h3f17_cfa3_786f_f108_bfb3_fdb2_4fb0_d0ef;
        state = 128'h0d8e_6d4a_c83c_5ebe_81f2_753a_dfc5_0490;

        #200;
        key = 128'hc05a_8896_34bf_0f18_05e5_300f_dd70_e5ad;
        state = 128'ha19c_0a2d_3ead_9545_c4ee_db04_c38c_3f33;

        #200;
        key = 128'h3009_8845_949e_1a5d_2a8c_931c_8104_346e;
        state = 128'h25c3_8c43_9209_3484_53e4_b2ad_c674_4a52;

        #200;
        key = 128'he4de_a1d2_026b_210c_5acd_2cec_91d6_dc4c;
        state = 128'h11ca_06b3_7bcf_90cc_c569_a1ac_7c4f_48c0;

        #200;
        key = 128'he3f3_73c6_545d_5ca6_dd9e_3ef4_d5f6_fd06;
        state = 128'h82d7_2fc6_b255_de54_8fec_d782_a146_1260;

        #200;
        key = 128'hd02c_2d50_c7e5_d881_877f_3046_df3b_4a37;
        state = 128'hcda6_f97b_d8a0_7afa_1a93_d38b_939e_5031;

        #200;
        key = 128'h53d9_d798_f946_4a82_965a_aba7_843d_9ff5;
        state = 128'hfc07_c846_92bb_a6e9_f783_4075_19e6_54f6;

        #200;
        key = 128'hd226_e05e_ac9d_9f02_4349_4293_876a_0f9c;
        state = 128'h3dfb_6def_0827_4084_785a_9736_0d13_c54f;

        #200;
        key = 128'h4b9d_ed20_0c84_9cb5_0b93_f480_1f0f_bad6;
        state = 128'h20de_6d19_b2ec_c1cb_c916_9557_5e49_b985;

        #200;
        key = 128'hedd5_0d40_b1d1_ff10_7e00_f55d_cde4_40eb;
        state = 128'hb692_5297_eea7_4459_768f_c541_16b9_d162;

        #200;
        key = 128'h16ea_4e19_89e0_b913_3ac8_5d25_459b_c0a5;
        state = 128'h497d_5f99_3f05_f9dd_2b9d_aeeb_eb36_c534;

        #200;
        key = 128'h5305_65ac_f7dd_3a20_01ec_c105_9cea_f97a;
        state = 128'h79fc_87c4_ae8c_eb90_a547_837b_b23a_e620;

        #200;
        key = 128'hc054_c4b4_b58b_101c_a03a_3e45_322e_4977;
        state = 128'hac6f_19fa_0d22_03b9_4d6c_6199_10b6_a5b6;

        #200;
        key = 128'ha3bc_0963_21f8_ce7e_169a_ad6f_b2f3_b6ea;
        state = 128'h7511_b1b0_f152_97bb_df38_818c_10df_089b;

        #200;
        key = 128'h6edb_f6e5_2402_6a30_5922_15b7_c74f_ad88;
        state = 128'h7098_8652_363b_1ffc_46e8_42e1_098d_ea69;

        #200;
        key = 128'h4a7e_0a67_2c44_b468_1a30_7eb2_c7f9_ff2d;
        state = 128'he740_9580_dacd_a2dc_2e6d_784c_011a_1984;

        #200;
        key = 128'h45d6_346f_3755_a759_05a8_1171_1191_52fc;
        state = 128'h2c76_8221_205c_247c_830c_2faa_eef3_e65f;

        #200;
        key = 128'haefb_4d13_b43f_9ccd_8a45_e065_bb06_c9e0;
        state = 128'h2e7d_9507_8e73_e22b_a1da_ffde_afa2_de65;

        #200;
        key = 128'h3c5f_1c98_aae3_fc28_d1d0_efd1_7bcf_dad8;
        state = 128'h9669_237d_be91_b402_f05a_2ad8_6c7b_27b3;

        #200;
        key = 128'hc427_62e7_f3f4_c0cb_3370_d235_8f21_891c;
        state = 128'h9d59_e2c8_6e85_af7b_039a_9a1d_e7d2_435d;

        #200;
        key = 128'hfde7_d489_fdad_dcb1_da00_87dd_8f4c_24a2;
        state = 128'h9b9b_5114_757a_593f_a566_6774_5df3_a7dd;

        #200;
        key = 128'ha06b_2021_dc1b_ced9_f71c_4806_6114_a1a0;
        state = 128'hc937_a06a_a93b_e3ec_108b_ecde_5997_15a5;

        #200;
        key = 128'h23fb_7980_f701_2a54_60a1_0394_dc8d_e23b;
        state = 128'hb4bd_60ad_de3d_d61a_b375_55ef_849a_9640;

        #200;
        key = 128'h2993_1838_438e_16bc_f794_8de3_a608_b0f5;
        state = 128'he2ad_5118_5130_b031_f572_b279_e668_0897;

        #200;
        key = 128'h7d35_eb3d_82b2_6b81_a861_beb3_9fd7_6c5f;
        state = 128'hd156_add6_a6bd_6e33_7595_9545_0984_f88d;

        #200;
        key = 128'h594e_a080_3e07_3f28_14fd_701b_04cc_b2b2;
        state = 128'he07e_2cc4_63e7_ba66_4e2f_c8c2_9f08_1e08;

        #200;
        key = 128'h67f6_38a7_74db_4e85_8858_2903_4129_3140;
        state = 128'h9e46_942e_26c8_1d52_e87a_e622_6628_1c88;

        #200;
        key = 128'h32a3_8d71_cc38_bf3d_c6c5_92b6_78ff_5253;
        state = 128'hf601_5e3b_a2b7_f012_3a10_3638_37d0_e2f6;

        #200;
        key = 128'h1504_37c6_4ac8_b668_bab0_eb85_3c36_9678;
        state = 128'h8cb8_2bdd_2ac8_4d9b_fe35_ff1d_fedb_54ba;

        #200;
        key = 128'h47c2_9ea0_e470_189a_cace_364a_d2af_b273;
        state = 128'h5cff_ef55_72f9_8e44_4d84_6f92_4c8c_f6c5;

        #200;
        key = 128'he061_cbeb_9c1b_4547_2389_d2b0_49fc_800b;
        state = 128'h7248_43aa_c6ac_bff2_cd6f_ac96_bcf2_29a2;

        #210 $finish;
    end 

endmodule
